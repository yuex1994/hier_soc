module oc8051__DOT__I__DOT__240(
__START__,
clk,
oc8051_ROM_rdata_0,
oc8051_ROM_rdata_1,
oc8051_ROM_rdata_2,
rst,
__ILA_oc8051_decode_of_I__DOT__240__,
__ILA_oc8051_valid__,
XRAM_addr0,
XRAM_data0,
XRAM_wen0,
ACC,
B,
DPH,
DPL,
IE,
IP,
P0,
P1,
P2,
P3,
PC,
PCON,
PSW,
SBUF,
SCON,
SP,
TCON,
TH0,
TH1,
TL0,
TL1,
TMOD,
XRAM_ADDR,
XRAM_DATA_IN,
XRAM_DATA_OUT,
oc8051_IRAM_data_0,
oc8051_IRAM_data_1,
oc8051_IRAM_data_2,
oc8051_IRAM_data_3,
oc8051_IRAM_data_4,
oc8051_IRAM_data_5,
oc8051_IRAM_data_6,
oc8051_IRAM_data_7,
oc8051_IRAM_data_8,
oc8051_IRAM_data_9,
oc8051_IRAM_data_10,
oc8051_IRAM_data_11,
oc8051_IRAM_data_12,
oc8051_IRAM_data_13,
oc8051_IRAM_data_14,
oc8051_IRAM_data_15,
oc8051_ROM_addr_0,
oc8051_ROM_addr_1,
oc8051_ROM_addr_2,
aes_address,
aes_length,
aes_key,
aes_counter,
aes_status,
__COUNTER_start__n1
);
input            __START__;
input            clk;
input      [7:0] oc8051_ROM_rdata_0;
input      [7:0] oc8051_ROM_rdata_1;
input      [7:0] oc8051_ROM_rdata_2;
input            rst;
output            __ILA_oc8051_decode_of_I__DOT__240__;
output            __ILA_oc8051_valid__;
output     [15:0] XRAM_addr0;
output      [7:0] XRAM_data0;
output            XRAM_wen0;
output reg      [7:0] ACC;
output reg      [7:0] B;
output reg      [7:0] DPH;
output reg      [7:0] DPL;
output reg      [7:0] IE;
output reg      [7:0] IP;
output reg      [7:0] P0;
output reg      [7:0] P1;
output reg      [7:0] P2;
output reg      [7:0] P3;
output reg     [15:0] PC;
output reg      [7:0] PCON;
output reg      [7:0] PSW;
output reg      [7:0] SBUF;
output reg      [7:0] SCON;
output reg      [7:0] SP;
output reg      [7:0] TCON;
output reg      [7:0] TH0;
output reg      [7:0] TH1;
output reg      [7:0] TL0;
output reg      [7:0] TL1;
output reg      [7:0] TMOD;
output reg     [15:0] XRAM_ADDR;
output reg      [7:0] XRAM_DATA_IN;
output reg      [7:0] XRAM_DATA_OUT;
output reg      [7:0] oc8051_IRAM_data_0;
output reg      [7:0] oc8051_IRAM_data_1;
output reg      [7:0] oc8051_IRAM_data_2;
output reg      [7:0] oc8051_IRAM_data_3;
output reg      [7:0] oc8051_IRAM_data_4;
output reg      [7:0] oc8051_IRAM_data_5;
output reg      [7:0] oc8051_IRAM_data_6;
output reg      [7:0] oc8051_IRAM_data_7;
output reg      [7:0] oc8051_IRAM_data_8;
output reg      [7:0] oc8051_IRAM_data_9;
output reg      [7:0] oc8051_IRAM_data_10;
output reg      [7:0] oc8051_IRAM_data_11;
output reg      [7:0] oc8051_IRAM_data_12;
output reg      [7:0] oc8051_IRAM_data_13;
output reg      [7:0] oc8051_IRAM_data_14;
output reg      [7:0] oc8051_IRAM_data_15;
output reg     [15:0] oc8051_ROM_addr_0;
output reg     [15:0] oc8051_ROM_addr_1;
output reg     [15:0] oc8051_ROM_addr_2;
output reg     [15:0] aes_address;
output reg     [15:0] aes_length;
output reg    [127:0] aes_key;
output reg    [127:0] aes_counter;
output reg      [1:0] aes_status;
output reg      [7:0] __COUNTER_start__n1;
(* keep *) wire      [7:0] ACC_randinit;
(* keep *) wire      [7:0] B_randinit;
(* keep *) wire      [7:0] DPH_randinit;
(* keep *) wire      [7:0] DPL_randinit;
(* keep *) wire      [7:0] IE_randinit;
(* keep *) wire      [7:0] IP_randinit;
(* keep *) wire      [7:0] P0_randinit;
(* keep *) wire      [7:0] P1_randinit;
(* keep *) wire      [7:0] P2_randinit;
(* keep *) wire      [7:0] P3_randinit;
(* keep *) wire      [7:0] PCON_randinit;
(* keep *) wire     [15:0] PC_randinit;
(* keep *) wire      [7:0] PSW_randinit;
(* keep *) wire      [7:0] SBUF_randinit;
(* keep *) wire      [7:0] SCON_randinit;
(* keep *) wire      [7:0] SP_randinit;
(* keep *) wire      [7:0] TCON_randinit;
(* keep *) wire      [7:0] TH0_randinit;
(* keep *) wire      [7:0] TH1_randinit;
(* keep *) wire      [7:0] TL0_randinit;
(* keep *) wire      [7:0] TL1_randinit;
(* keep *) wire      [7:0] TMOD_randinit;
(* keep *) wire     [15:0] XRAM_ADDR_randinit;
(* keep *) wire      [7:0] XRAM_DATA_IN_randinit;
(* keep *) wire      [7:0] XRAM_DATA_OUT_randinit;
wire     [15:0] XRAM_addr0;
wire      [7:0] XRAM_data0;
wire            XRAM_wen0;
wire            __ILA_oc8051_decode_of_I__DOT__240__;
wire            __ILA_oc8051_valid__;
wire            __START__;
(* keep *) wire     [15:0] aes_address_randinit;
(* keep *) wire    [127:0] aes_counter_randinit;
(* keep *) wire    [127:0] aes_key_randinit;
(* keep *) wire     [15:0] aes_length_randinit;
(* keep *) wire      [1:0] aes_status_randinit;
wire            clk;
wire            n0____DOLLAR__167758;
wire     [15:0] n1000____DOLLAR__2450;
wire            n1001____DOLLAR__2456;
wire            n1002____DOLLAR__2460;
wire            n1003____DOLLAR__2462;
wire            n1004____DOLLAR__2468;
wire            n1005____DOLLAR__2472;
wire      [4:0] n1006____DOLLAR__2474;
wire      [7:0] n1007____DOLLAR__2482;
wire      [7:0] n1008____DOLLAR__2484;
wire      [7:0] n1009____DOLLAR__2488;
wire            n100____DOLLAR__469;
wire      [7:0] n1010____DOLLAR__2489;
wire            n1011____DOLLAR__2490;
wire            n1012____DOLLAR__2494;
wire      [3:0] n1013____DOLLAR__178417;
wire            n1014____DOLLAR__178498;
wire            n1015____DOLLAR__178493;
wire            n1016____DOLLAR__178488;
wire            n1017____DOLLAR__178483;
wire            n1018____DOLLAR__178478;
wire            n1019____DOLLAR__178473;
wire            n101____DOLLAR__473;
wire            n1020____DOLLAR__178468;
wire            n1021____DOLLAR__178463;
wire            n1022____DOLLAR__178458;
wire            n1023____DOLLAR__178453;
wire            n1024____DOLLAR__178448;
wire            n1025____DOLLAR__178443;
wire            n1026____DOLLAR__178438;
wire            n1027____DOLLAR__178433;
wire            n1028____DOLLAR__178428;
wire            n1029____DOLLAR__178423;
wire            n102____DOLLAR__477;
wire      [7:0] n1030____DOLLAR__178425;
wire      [7:0] n1031____DOLLAR__178430;
wire      [7:0] n1032____DOLLAR__178435;
wire      [7:0] n1033____DOLLAR__178440;
wire      [7:0] n1034____DOLLAR__178445;
wire      [7:0] n1035____DOLLAR__178450;
wire      [7:0] n1036____DOLLAR__178455;
wire      [7:0] n1037____DOLLAR__178460;
wire      [7:0] n1038____DOLLAR__178465;
wire      [7:0] n1039____DOLLAR__178470;
wire            n103____DOLLAR__481;
wire      [7:0] n1040____DOLLAR__178475;
wire      [7:0] n1041____DOLLAR__178480;
wire      [7:0] n1042____DOLLAR__178485;
wire      [7:0] n1043____DOLLAR__178490;
wire      [7:0] n1044____DOLLAR__178495;
wire      [7:0] n1045____DOLLAR__178500;
wire            n1046____DOLLAR__2500;
wire            n1047____DOLLAR__2504;
wire            n1048____DOLLAR__2508;
wire            n1049____DOLLAR__2512;
wire            n104____DOLLAR__485;
wire            n1050____DOLLAR__2516;
wire            n1051____DOLLAR__2520;
wire            n1052____DOLLAR__2524;
wire            n1053____DOLLAR__2528;
wire            n1054____DOLLAR__2532;
wire            n1055____DOLLAR__2536;
wire            n1056____DOLLAR__2540;
wire            n1057____DOLLAR__2544;
wire            n1058____DOLLAR__2548;
wire            n1059____DOLLAR__2552;
wire            n105____DOLLAR__489;
wire            n1060____DOLLAR__2556;
wire            n1061____DOLLAR__2560;
wire            n1062____DOLLAR__2564;
wire            n1063____DOLLAR__2568;
wire            n1064____DOLLAR__2572;
wire            n1065____DOLLAR__2576;
wire            n1066____DOLLAR__2580;
wire      [7:0] n1067____DOLLAR__2584;
wire      [7:0] n1068____DOLLAR__2585;
wire      [7:0] n1069____DOLLAR__2586;
wire            n106____DOLLAR__493;
wire      [7:0] n1070____DOLLAR__2587;
wire      [7:0] n1071____DOLLAR__2588;
wire      [7:0] n1072____DOLLAR__2589;
wire      [7:0] n1073____DOLLAR__2590;
wire      [7:0] n1074____DOLLAR__2591;
wire      [7:0] n1075____DOLLAR__2592;
wire      [7:0] n1076____DOLLAR__2593;
wire      [7:0] n1077____DOLLAR__2594;
wire      [7:0] n1078____DOLLAR__2595;
wire      [7:0] n1079____DOLLAR__2596;
wire            n107____DOLLAR__497;
wire      [7:0] n1080____DOLLAR__2597;
wire      [7:0] n1081____DOLLAR__2598;
wire      [7:0] n1082____DOLLAR__2599;
wire      [7:0] n1083____DOLLAR__2600;
wire      [7:0] n1084____DOLLAR__2601;
wire      [7:0] n1085____DOLLAR__2602;
wire      [7:0] n1086____DOLLAR__2603;
wire      [7:0] n1087____DOLLAR__2604;
wire      [7:0] n1088____DOLLAR__2605;
wire            n1089____DOLLAR__2606;
wire            n108____DOLLAR__501;
wire            n1090____DOLLAR__2608;
wire     [15:0] n1091____DOLLAR__2612;
wire     [15:0] n1092____DOLLAR__2618;
wire     [15:0] n1093____DOLLAR__2620;
wire     [15:0] n1094____DOLLAR__2623;
wire     [15:0] n1095____DOLLAR__2624;
wire            n1096____DOLLAR__2629;
wire            n1097____DOLLAR__2633;
wire            n1098____DOLLAR__2637;
wire            n1099____DOLLAR__2641;
wire            n109____DOLLAR__505;
wire            n10____DOLLAR__109;
wire            n1100____DOLLAR__2645;
wire            n1101____DOLLAR__2649;
wire            n1102____DOLLAR__2653;
wire            n1103____DOLLAR__2657;
wire            n1104____DOLLAR__2661;
wire            n1105____DOLLAR__2665;
wire            n1106____DOLLAR__2669;
wire            n1107____DOLLAR__2673;
wire            n1108____DOLLAR__2677;
wire            n1109____DOLLAR__2681;
wire            n110____DOLLAR__509;
wire            n1110____DOLLAR__2685;
wire            n1111____DOLLAR__2689;
wire            n1112____DOLLAR__2693;
wire            n1113____DOLLAR__2697;
wire            n1114____DOLLAR__2701;
wire            n1115____DOLLAR__2705;
wire            n1116____DOLLAR__2709;
wire            n1117____DOLLAR__2713;
wire            n1118____DOLLAR__2717;
wire            n1119____DOLLAR__2721;
wire            n111____DOLLAR__513;
wire            n1120____DOLLAR__2725;
wire            n1121____DOLLAR__2729;
wire            n1122____DOLLAR__2733;
wire            n1123____DOLLAR__2737;
wire            n1124____DOLLAR__2741;
wire            n1125____DOLLAR__2745;
wire            n1126____DOLLAR__2749;
wire            n1127____DOLLAR__2753;
wire            n1128____DOLLAR__2757;
wire            n1129____DOLLAR__2761;
wire            n112____DOLLAR__517;
wire            n1130____DOLLAR__2765;
wire            n1131____DOLLAR__2769;
wire            n1132____DOLLAR__2773;
wire            n1133____DOLLAR__2777;
wire            n1134____DOLLAR__2781;
wire            n1135____DOLLAR__2785;
wire            n1136____DOLLAR__2789;
wire            n1137____DOLLAR__2793;
wire            n1138____DOLLAR__2797;
wire            n1139____DOLLAR__2801;
wire            n113____DOLLAR__521;
wire            n1140____DOLLAR__2805;
wire            n1141____DOLLAR__2809;
wire            n1142____DOLLAR__2813;
wire            n1143____DOLLAR__2817;
wire            n1144____DOLLAR__2821;
wire            n1145____DOLLAR__2825;
wire            n1146____DOLLAR__2829;
wire            n1147____DOLLAR__2833;
wire            n1148____DOLLAR__2837;
wire            n1149____DOLLAR__2841;
wire            n114____DOLLAR__525;
wire            n1150____DOLLAR__2845;
wire            n1151____DOLLAR__2849;
wire            n1152____DOLLAR__2853;
wire            n1153____DOLLAR__2857;
wire            n1154____DOLLAR__2861;
wire            n1155____DOLLAR__2865;
wire            n1156____DOLLAR__2869;
wire            n1157____DOLLAR__2873;
wire            n1158____DOLLAR__2875;
wire            n1159____DOLLAR__2876;
wire            n115____DOLLAR__529;
wire            n1160____DOLLAR__2877;
wire            n1161____DOLLAR__2878;
wire            n1162____DOLLAR__2879;
wire            n1163____DOLLAR__2880;
wire            n1164____DOLLAR__2881;
wire            n1165____DOLLAR__2882;
wire            n1166____DOLLAR__2883;
wire            n1167____DOLLAR__2884;
wire            n1168____DOLLAR__2885;
wire            n1169____DOLLAR__2886;
wire            n116____DOLLAR__533;
wire            n1170____DOLLAR__2887;
wire            n1171____DOLLAR__2888;
wire            n1172____DOLLAR__2889;
wire            n1173____DOLLAR__2890;
wire            n1174____DOLLAR__2891;
wire            n1175____DOLLAR__2892;
wire            n1176____DOLLAR__2893;
wire            n1177____DOLLAR__2894;
wire            n1178____DOLLAR__2895;
wire            n1179____DOLLAR__2896;
wire            n117____DOLLAR__537;
wire            n1180____DOLLAR__2897;
wire            n1181____DOLLAR__2898;
wire            n1182____DOLLAR__2899;
wire            n1183____DOLLAR__2900;
wire            n1184____DOLLAR__2901;
wire            n1185____DOLLAR__2902;
wire            n1186____DOLLAR__2903;
wire            n1187____DOLLAR__2904;
wire            n1188____DOLLAR__2905;
wire            n1189____DOLLAR__2906;
wire            n118____DOLLAR__541;
wire            n1190____DOLLAR__2907;
wire            n1191____DOLLAR__2908;
wire            n1192____DOLLAR__2909;
wire            n1193____DOLLAR__2910;
wire            n1194____DOLLAR__2911;
wire            n1195____DOLLAR__2912;
wire            n1196____DOLLAR__2913;
wire            n1197____DOLLAR__2914;
wire            n1198____DOLLAR__2915;
wire            n1199____DOLLAR__2916;
wire            n119____DOLLAR__545;
wire            n11____DOLLAR__113;
wire            n1200____DOLLAR__2917;
wire            n1201____DOLLAR__2918;
wire            n1202____DOLLAR__2919;
wire            n1203____DOLLAR__2920;
wire            n1204____DOLLAR__2921;
wire            n1205____DOLLAR__2922;
wire            n1206____DOLLAR__2923;
wire            n1207____DOLLAR__2924;
wire            n1208____DOLLAR__2925;
wire            n1209____DOLLAR__2926;
wire            n120____DOLLAR__549;
wire            n1210____DOLLAR__2927;
wire            n1211____DOLLAR__2928;
wire            n1212____DOLLAR__2929;
wire            n1213____DOLLAR__2930;
wire            n1214____DOLLAR__2931;
wire            n1215____DOLLAR__2932;
wire            n1216____DOLLAR__2933;
wire            n1217____DOLLAR__2934;
wire            n1218____DOLLAR__2935;
wire     [15:0] n1219____DOLLAR__2938;
wire            n121____DOLLAR__553;
wire            n1220____DOLLAR__2943;
wire            n1221____DOLLAR__2947;
wire            n1222____DOLLAR__2949;
wire     [15:0] n1223____DOLLAR__2964;
wire            n1224____DOLLAR__2970;
wire            n1225____DOLLAR__2974;
wire            n1226____DOLLAR__2976;
wire     [15:0] n1227____DOLLAR__2979;
wire      [4:0] n1228____DOLLAR__2980;
wire      [7:0] n1229____DOLLAR__2988;
wire            n122____DOLLAR__557;
wire     [15:0] n1230____DOLLAR__2999;
wire            n1231____DOLLAR__3005;
wire            n1232____DOLLAR__3009;
wire            n1233____DOLLAR__3013;
wire            n1234____DOLLAR__3017;
wire            n1235____DOLLAR__3021;
wire            n1236____DOLLAR__3025;
wire            n1237____DOLLAR__3029;
wire            n1238____DOLLAR__3033;
wire            n1239____DOLLAR__3037;
wire            n123____DOLLAR__561;
wire            n1240____DOLLAR__3041;
wire            n1241____DOLLAR__3045;
wire            n1242____DOLLAR__3049;
wire            n1243____DOLLAR__3053;
wire            n1244____DOLLAR__3057;
wire            n1245____DOLLAR__3061;
wire            n1246____DOLLAR__3065;
wire            n1247____DOLLAR__3069;
wire            n1248____DOLLAR__3073;
wire            n1249____DOLLAR__3077;
wire            n124____DOLLAR__565;
wire            n1250____DOLLAR__3081;
wire            n1251____DOLLAR__3085;
wire            n1252____DOLLAR__3089;
wire            n1253____DOLLAR__3093;
wire            n1254____DOLLAR__3097;
wire            n1255____DOLLAR__3101;
wire            n1256____DOLLAR__3105;
wire            n1257____DOLLAR__3109;
wire            n1258____DOLLAR__3113;
wire            n1259____DOLLAR__3117;
wire            n125____DOLLAR__569;
wire            n1260____DOLLAR__3121;
wire            n1261____DOLLAR__3125;
wire            n1262____DOLLAR__3129;
wire            n1263____DOLLAR__3133;
wire            n1264____DOLLAR__3137;
wire            n1265____DOLLAR__3141;
wire            n1266____DOLLAR__3145;
wire            n1267____DOLLAR__3149;
wire            n1268____DOLLAR__3153;
wire            n1269____DOLLAR__3157;
wire            n126____DOLLAR__573;
wire            n1270____DOLLAR__3161;
wire            n1271____DOLLAR__3165;
wire            n1272____DOLLAR__3169;
wire            n1273____DOLLAR__3173;
wire            n1274____DOLLAR__3177;
wire            n1275____DOLLAR__3181;
wire            n1276____DOLLAR__3185;
wire            n1277____DOLLAR__3189;
wire            n1278____DOLLAR__3193;
wire            n1279____DOLLAR__3197;
wire            n127____DOLLAR__577;
wire            n1280____DOLLAR__3201;
wire            n1281____DOLLAR__3205;
wire            n1282____DOLLAR__3209;
wire            n1283____DOLLAR__3213;
wire            n1284____DOLLAR__3217;
wire            n1285____DOLLAR__3221;
wire            n1286____DOLLAR__3225;
wire            n1287____DOLLAR__3229;
wire            n1288____DOLLAR__3233;
wire            n1289____DOLLAR__3237;
wire            n128____DOLLAR__581;
wire            n1290____DOLLAR__3241;
wire            n1291____DOLLAR__3245;
wire            n1292____DOLLAR__3249;
wire            n1293____DOLLAR__3253;
wire            n1294____DOLLAR__3257;
wire            n1295____DOLLAR__3261;
wire            n1296____DOLLAR__3265;
wire            n1297____DOLLAR__3269;
wire            n1298____DOLLAR__3273;
wire            n1299____DOLLAR__3277;
wire            n129____DOLLAR__585;
wire            n12____DOLLAR__117;
wire            n1300____DOLLAR__3281;
wire            n1301____DOLLAR__3285;
wire            n1302____DOLLAR__3289;
wire            n1303____DOLLAR__3293;
wire            n1304____DOLLAR__3297;
wire            n1305____DOLLAR__3301;
wire            n1306____DOLLAR__3305;
wire            n1307____DOLLAR__3309;
wire            n1308____DOLLAR__3313;
wire            n1309____DOLLAR__3317;
wire            n130____DOLLAR__589;
wire            n1310____DOLLAR__3321;
wire            n1311____DOLLAR__3325;
wire            n1312____DOLLAR__3329;
wire            n1313____DOLLAR__3333;
wire            n1314____DOLLAR__3337;
wire            n1315____DOLLAR__3341;
wire            n1316____DOLLAR__3345;
wire            n1317____DOLLAR__3349;
wire            n1318____DOLLAR__3353;
wire            n1319____DOLLAR__3357;
wire            n131____DOLLAR__593;
wire            n1320____DOLLAR__3361;
wire            n1321____DOLLAR__3365;
wire            n1322____DOLLAR__3369;
wire            n1323____DOLLAR__3373;
wire            n1324____DOLLAR__3377;
wire            n1325____DOLLAR__3381;
wire            n1326____DOLLAR__3385;
wire            n1327____DOLLAR__3389;
wire            n1328____DOLLAR__3393;
wire            n1329____DOLLAR__3397;
wire            n132____DOLLAR__597;
wire            n1330____DOLLAR__3401;
wire            n1331____DOLLAR__3405;
wire            n1332____DOLLAR__3409;
wire            n1333____DOLLAR__3413;
wire            n1334____DOLLAR__3417;
wire            n1335____DOLLAR__3421;
wire            n1336____DOLLAR__3425;
wire            n1337____DOLLAR__3429;
wire            n1338____DOLLAR__3433;
wire            n1339____DOLLAR__3437;
wire            n133____DOLLAR__601;
wire            n1340____DOLLAR__3441;
wire            n1341____DOLLAR__3445;
wire            n1342____DOLLAR__3449;
wire            n1343____DOLLAR__3453;
wire            n1344____DOLLAR__3457;
wire            n1345____DOLLAR__3461;
wire            n1346____DOLLAR__3465;
wire            n1347____DOLLAR__3469;
wire            n1348____DOLLAR__3473;
wire            n1349____DOLLAR__3477;
wire            n134____DOLLAR__605;
wire            n1350____DOLLAR__3481;
wire            n1351____DOLLAR__3485;
wire            n1352____DOLLAR__3489;
wire            n1353____DOLLAR__3493;
wire            n1354____DOLLAR__3497;
wire            n1355____DOLLAR__3501;
wire            n1356____DOLLAR__3505;
wire            n1357____DOLLAR__3509;
wire            n1358____DOLLAR__3513;
wire            n1359____DOLLAR__3517;
wire            n135____DOLLAR__609;
wire            n1360____DOLLAR__3521;
wire            n1361____DOLLAR__3525;
wire            n1362____DOLLAR__3529;
wire            n1363____DOLLAR__3533;
wire            n1364____DOLLAR__3537;
wire            n1365____DOLLAR__3541;
wire            n1366____DOLLAR__3545;
wire            n1367____DOLLAR__3549;
wire            n1368____DOLLAR__3553;
wire            n1369____DOLLAR__3555;
wire            n136____DOLLAR__613;
wire            n1370____DOLLAR__3556;
wire            n1371____DOLLAR__3557;
wire            n1372____DOLLAR__3558;
wire            n1373____DOLLAR__3559;
wire            n1374____DOLLAR__3560;
wire            n1375____DOLLAR__3561;
wire            n1376____DOLLAR__3562;
wire            n1377____DOLLAR__3563;
wire            n1378____DOLLAR__3564;
wire            n1379____DOLLAR__3565;
wire            n137____DOLLAR__617;
wire            n1380____DOLLAR__3566;
wire            n1381____DOLLAR__3567;
wire            n1382____DOLLAR__3568;
wire            n1383____DOLLAR__3569;
wire            n1384____DOLLAR__3570;
wire            n1385____DOLLAR__3571;
wire            n1386____DOLLAR__3572;
wire            n1387____DOLLAR__3573;
wire            n1388____DOLLAR__3574;
wire            n1389____DOLLAR__3575;
wire            n138____DOLLAR__621;
wire            n1390____DOLLAR__3576;
wire            n1391____DOLLAR__3577;
wire            n1392____DOLLAR__3578;
wire            n1393____DOLLAR__3579;
wire            n1394____DOLLAR__3580;
wire            n1395____DOLLAR__3581;
wire            n1396____DOLLAR__3582;
wire            n1397____DOLLAR__3583;
wire            n1398____DOLLAR__3584;
wire            n1399____DOLLAR__3585;
wire            n139____DOLLAR__625;
wire            n13____DOLLAR__121;
wire            n1400____DOLLAR__3586;
wire            n1401____DOLLAR__3587;
wire            n1402____DOLLAR__3588;
wire            n1403____DOLLAR__3589;
wire            n1404____DOLLAR__3590;
wire            n1405____DOLLAR__3591;
wire            n1406____DOLLAR__3592;
wire            n1407____DOLLAR__3593;
wire            n1408____DOLLAR__3594;
wire            n1409____DOLLAR__3595;
wire            n140____DOLLAR__629;
wire            n1410____DOLLAR__3596;
wire            n1411____DOLLAR__3597;
wire            n1412____DOLLAR__3598;
wire            n1413____DOLLAR__3599;
wire            n1414____DOLLAR__3600;
wire            n1415____DOLLAR__3601;
wire            n1416____DOLLAR__3602;
wire            n1417____DOLLAR__3603;
wire            n1418____DOLLAR__3604;
wire            n1419____DOLLAR__3605;
wire            n141____DOLLAR__633;
wire            n1420____DOLLAR__3606;
wire            n1421____DOLLAR__3607;
wire            n1422____DOLLAR__3608;
wire            n1423____DOLLAR__3609;
wire            n1424____DOLLAR__3610;
wire            n1425____DOLLAR__3611;
wire            n1426____DOLLAR__3612;
wire            n1427____DOLLAR__3613;
wire            n1428____DOLLAR__3614;
wire            n1429____DOLLAR__3615;
wire            n142____DOLLAR__637;
wire            n1430____DOLLAR__3616;
wire            n1431____DOLLAR__3617;
wire            n1432____DOLLAR__3618;
wire            n1433____DOLLAR__3619;
wire            n1434____DOLLAR__3620;
wire            n1435____DOLLAR__3621;
wire            n1436____DOLLAR__3622;
wire            n1437____DOLLAR__3623;
wire            n1438____DOLLAR__3624;
wire            n1439____DOLLAR__3625;
wire            n143____DOLLAR__641;
wire            n1440____DOLLAR__3626;
wire            n1441____DOLLAR__3627;
wire            n1442____DOLLAR__3628;
wire            n1443____DOLLAR__3629;
wire            n1444____DOLLAR__3630;
wire            n1445____DOLLAR__3631;
wire            n1446____DOLLAR__3632;
wire            n1447____DOLLAR__3633;
wire            n1448____DOLLAR__3634;
wire            n1449____DOLLAR__3635;
wire            n144____DOLLAR__645;
wire            n1450____DOLLAR__3636;
wire            n1451____DOLLAR__3637;
wire            n1452____DOLLAR__3638;
wire            n1453____DOLLAR__3639;
wire            n1454____DOLLAR__3640;
wire            n1455____DOLLAR__3641;
wire            n1456____DOLLAR__3642;
wire            n1457____DOLLAR__3643;
wire            n1458____DOLLAR__3644;
wire            n1459____DOLLAR__3645;
wire            n145____DOLLAR__649;
wire            n1460____DOLLAR__3646;
wire            n1461____DOLLAR__3647;
wire            n1462____DOLLAR__3648;
wire            n1463____DOLLAR__3649;
wire            n1464____DOLLAR__3650;
wire            n1465____DOLLAR__3651;
wire            n1466____DOLLAR__3652;
wire            n1467____DOLLAR__3653;
wire            n1468____DOLLAR__3654;
wire            n1469____DOLLAR__3655;
wire            n146____DOLLAR__653;
wire            n1470____DOLLAR__3656;
wire            n1471____DOLLAR__3657;
wire            n1472____DOLLAR__3658;
wire            n1473____DOLLAR__3659;
wire            n1474____DOLLAR__3660;
wire            n1475____DOLLAR__3661;
wire            n1476____DOLLAR__3662;
wire            n1477____DOLLAR__3663;
wire            n1478____DOLLAR__3664;
wire            n1479____DOLLAR__3665;
wire            n147____DOLLAR__657;
wire            n1480____DOLLAR__3666;
wire            n1481____DOLLAR__3667;
wire            n1482____DOLLAR__3668;
wire            n1483____DOLLAR__3669;
wire            n1484____DOLLAR__3670;
wire            n1485____DOLLAR__3671;
wire            n1486____DOLLAR__3672;
wire            n1487____DOLLAR__3673;
wire            n1488____DOLLAR__3674;
wire            n1489____DOLLAR__3675;
wire            n148____DOLLAR__661;
wire            n1490____DOLLAR__3676;
wire            n1491____DOLLAR__3677;
wire            n1492____DOLLAR__3678;
wire            n1493____DOLLAR__3679;
wire            n1494____DOLLAR__3680;
wire            n1495____DOLLAR__3681;
wire            n1496____DOLLAR__3682;
wire            n1497____DOLLAR__3683;
wire            n1498____DOLLAR__3684;
wire            n1499____DOLLAR__3685;
wire            n149____DOLLAR__665;
wire            n14____DOLLAR__125;
wire            n1500____DOLLAR__3686;
wire            n1501____DOLLAR__3687;
wire            n1502____DOLLAR__3688;
wire            n1503____DOLLAR__3689;
wire            n1504____DOLLAR__3690;
wire            n1505____DOLLAR__3691;
wire     [15:0] n1506____DOLLAR__3694;
wire     [15:0] n1507____DOLLAR__3695;
wire     [15:0] n1508____DOLLAR__3696;
wire     [15:0] n1509____DOLLAR__3697;
wire            n150____DOLLAR__669;
wire     [15:0] n1510____DOLLAR__3698;
wire     [15:0] n1511____DOLLAR__3699;
wire     [15:0] n1512____DOLLAR__3700;
wire     [15:0] n1513____DOLLAR__3701;
wire            n1514____DOLLAR__3706;
wire            n1515____DOLLAR__3710;
wire            n1516____DOLLAR__3714;
wire            n1517____DOLLAR__3718;
wire            n1518____DOLLAR__3722;
wire            n1519____DOLLAR__3726;
wire            n151____DOLLAR__673;
wire            n1520____DOLLAR__3730;
wire            n1521____DOLLAR__3734;
wire            n1522____DOLLAR__3738;
wire            n1523____DOLLAR__3742;
wire            n1524____DOLLAR__3746;
wire            n1525____DOLLAR__3750;
wire            n1526____DOLLAR__3754;
wire            n1527____DOLLAR__3758;
wire            n1528____DOLLAR__3762;
wire            n1529____DOLLAR__3766;
wire            n152____DOLLAR__677;
wire            n1530____DOLLAR__3770;
wire            n1531____DOLLAR__3774;
wire            n1532____DOLLAR__3778;
wire            n1533____DOLLAR__3782;
wire            n1534____DOLLAR__3786;
wire            n1535____DOLLAR__3790;
wire            n1536____DOLLAR__3794;
wire            n1537____DOLLAR__3798;
wire            n1538____DOLLAR__3802;
wire            n1539____DOLLAR__3806;
wire            n153____DOLLAR__681;
wire            n1540____DOLLAR__3810;
wire            n1541____DOLLAR__3814;
wire            n1542____DOLLAR__3818;
wire            n1543____DOLLAR__3822;
wire            n1544____DOLLAR__3826;
wire            n1545____DOLLAR__3830;
wire            n1546____DOLLAR__3834;
wire            n1547____DOLLAR__3838;
wire            n1548____DOLLAR__3842;
wire            n1549____DOLLAR__3846;
wire            n154____DOLLAR__685;
wire            n1550____DOLLAR__3850;
wire            n1551____DOLLAR__3854;
wire            n1552____DOLLAR__3858;
wire            n1553____DOLLAR__3862;
wire            n1554____DOLLAR__3866;
wire            n1555____DOLLAR__3870;
wire            n1556____DOLLAR__3874;
wire            n1557____DOLLAR__3878;
wire            n1558____DOLLAR__3882;
wire            n1559____DOLLAR__3886;
wire            n155____DOLLAR__689;
wire            n1560____DOLLAR__3890;
wire            n1561____DOLLAR__3894;
wire            n1562____DOLLAR__3898;
wire            n1563____DOLLAR__3902;
wire            n1564____DOLLAR__3906;
wire            n1565____DOLLAR__3910;
wire            n1566____DOLLAR__3914;
wire            n1567____DOLLAR__3918;
wire            n1568____DOLLAR__3922;
wire            n1569____DOLLAR__3926;
wire            n156____DOLLAR__693;
wire            n1570____DOLLAR__3930;
wire            n1571____DOLLAR__3934;
wire            n1572____DOLLAR__3938;
wire            n1573____DOLLAR__3942;
wire            n1574____DOLLAR__3946;
wire            n1575____DOLLAR__3950;
wire            n1576____DOLLAR__3954;
wire            n1577____DOLLAR__3958;
wire            n1578____DOLLAR__3962;
wire            n1579____DOLLAR__3966;
wire            n157____DOLLAR__697;
wire            n1580____DOLLAR__3970;
wire            n1581____DOLLAR__3974;
wire            n1582____DOLLAR__3978;
wire            n1583____DOLLAR__3982;
wire            n1584____DOLLAR__3986;
wire            n1585____DOLLAR__3990;
wire            n1586____DOLLAR__3994;
wire            n1587____DOLLAR__3998;
wire            n1588____DOLLAR__4002;
wire            n1589____DOLLAR__4006;
wire            n158____DOLLAR__701;
wire            n1590____DOLLAR__4010;
wire            n1591____DOLLAR__4014;
wire            n1592____DOLLAR__4018;
wire            n1593____DOLLAR__4022;
wire            n1594____DOLLAR__4026;
wire            n1595____DOLLAR__4030;
wire            n1596____DOLLAR__4034;
wire            n1597____DOLLAR__4038;
wire            n1598____DOLLAR__4042;
wire            n1599____DOLLAR__4046;
wire            n159____DOLLAR__705;
wire            n15____DOLLAR__129;
wire            n1600____DOLLAR__4050;
wire            n1601____DOLLAR__4054;
wire            n1602____DOLLAR__4058;
wire            n1603____DOLLAR__4062;
wire            n1604____DOLLAR__4066;
wire            n1605____DOLLAR__4070;
wire            n1606____DOLLAR__4074;
wire            n1607____DOLLAR__4078;
wire            n1608____DOLLAR__4082;
wire            n1609____DOLLAR__4086;
wire            n160____DOLLAR__709;
wire            n1610____DOLLAR__4090;
wire            n1611____DOLLAR__4094;
wire            n1612____DOLLAR__4098;
wire            n1613____DOLLAR__4102;
wire            n1614____DOLLAR__4106;
wire            n1615____DOLLAR__4110;
wire            n1616____DOLLAR__4114;
wire            n1617____DOLLAR__4118;
wire            n1618____DOLLAR__4122;
wire            n1619____DOLLAR__4126;
wire            n161____DOLLAR__713;
wire            n1620____DOLLAR__4130;
wire            n1621____DOLLAR__4134;
wire            n1622____DOLLAR__4138;
wire            n1623____DOLLAR__4142;
wire            n1624____DOLLAR__4146;
wire            n1625____DOLLAR__4150;
wire            n1626____DOLLAR__4154;
wire            n1627____DOLLAR__4158;
wire            n1628____DOLLAR__4162;
wire            n1629____DOLLAR__4166;
wire            n162____DOLLAR__717;
wire            n1630____DOLLAR__4170;
wire            n1631____DOLLAR__4174;
wire            n1632____DOLLAR__4178;
wire            n1633____DOLLAR__4182;
wire            n1634____DOLLAR__4186;
wire            n1635____DOLLAR__4190;
wire            n1636____DOLLAR__4194;
wire            n1637____DOLLAR__4198;
wire            n1638____DOLLAR__4202;
wire            n1639____DOLLAR__4206;
wire            n163____DOLLAR__721;
wire            n1640____DOLLAR__4210;
wire            n1641____DOLLAR__4214;
wire            n1642____DOLLAR__4218;
wire            n1643____DOLLAR__4222;
wire            n1644____DOLLAR__4226;
wire            n1645____DOLLAR__4230;
wire            n1646____DOLLAR__4234;
wire            n1647____DOLLAR__4238;
wire            n1648____DOLLAR__4242;
wire            n1649____DOLLAR__4246;
wire            n164____DOLLAR__725;
wire            n1650____DOLLAR__4250;
wire            n1651____DOLLAR__4254;
wire            n1652____DOLLAR__4258;
wire            n1653____DOLLAR__4262;
wire            n1654____DOLLAR__4266;
wire            n1655____DOLLAR__4270;
wire            n1656____DOLLAR__4274;
wire            n1657____DOLLAR__4278;
wire            n1658____DOLLAR__4282;
wire            n1659____DOLLAR__4286;
wire            n165____DOLLAR__729;
wire            n1660____DOLLAR__4290;
wire            n1661____DOLLAR__4294;
wire            n1662____DOLLAR__4298;
wire            n1663____DOLLAR__4302;
wire            n1664____DOLLAR__4306;
wire            n1665____DOLLAR__4310;
wire            n1666____DOLLAR__4314;
wire            n1667____DOLLAR__4318;
wire            n1668____DOLLAR__4322;
wire            n1669____DOLLAR__4326;
wire            n166____DOLLAR__733;
wire            n1670____DOLLAR__4330;
wire            n1671____DOLLAR__4334;
wire            n1672____DOLLAR__4338;
wire            n1673____DOLLAR__4342;
wire            n1674____DOLLAR__4346;
wire            n1675____DOLLAR__4350;
wire            n1676____DOLLAR__4354;
wire            n1677____DOLLAR__4358;
wire            n1678____DOLLAR__4362;
wire            n1679____DOLLAR__4366;
wire            n167____DOLLAR__737;
wire            n1680____DOLLAR__4370;
wire            n1681____DOLLAR__4374;
wire            n1682____DOLLAR__4378;
wire            n1683____DOLLAR__4382;
wire            n1684____DOLLAR__4386;
wire            n1685____DOLLAR__4390;
wire            n1686____DOLLAR__4394;
wire            n1687____DOLLAR__4398;
wire            n1688____DOLLAR__4402;
wire            n1689____DOLLAR__4406;
wire            n168____DOLLAR__741;
wire            n1690____DOLLAR__4410;
wire            n1691____DOLLAR__4414;
wire            n1692____DOLLAR__4418;
wire            n1693____DOLLAR__4422;
wire            n1694____DOLLAR__4426;
wire            n1695____DOLLAR__4430;
wire            n1696____DOLLAR__4434;
wire            n1697____DOLLAR__4438;
wire            n1698____DOLLAR__4442;
wire            n1699____DOLLAR__4446;
wire            n169____DOLLAR__745;
wire            n16____DOLLAR__133;
wire            n1700____DOLLAR__4450;
wire            n1701____DOLLAR__4454;
wire            n1702____DOLLAR__4458;
wire            n1703____DOLLAR__4462;
wire            n1704____DOLLAR__4466;
wire            n1705____DOLLAR__4470;
wire            n1706____DOLLAR__4474;
wire            n1707____DOLLAR__4478;
wire            n1708____DOLLAR__4482;
wire            n1709____DOLLAR__4486;
wire            n170____DOLLAR__749;
wire            n1710____DOLLAR__4490;
wire            n1711____DOLLAR__4494;
wire            n1712____DOLLAR__4498;
wire            n1713____DOLLAR__4502;
wire            n1714____DOLLAR__4506;
wire            n1715____DOLLAR__4510;
wire            n1716____DOLLAR__4514;
wire            n1717____DOLLAR__4518;
wire            n1718____DOLLAR__4522;
wire            n1719____DOLLAR__4526;
wire            n171____DOLLAR__753;
wire            n1720____DOLLAR__4530;
wire            n1721____DOLLAR__4534;
wire            n1722____DOLLAR__4538;
wire            n1723____DOLLAR__4542;
wire            n1724____DOLLAR__4546;
wire            n1725____DOLLAR__4550;
wire            n1726____DOLLAR__4554;
wire            n1727____DOLLAR__4558;
wire            n1728____DOLLAR__4562;
wire            n1729____DOLLAR__4566;
wire            n172____DOLLAR__757;
wire            n1730____DOLLAR__4570;
wire            n1731____DOLLAR__4574;
wire            n1732____DOLLAR__4578;
wire            n1733____DOLLAR__4582;
wire            n1734____DOLLAR__4584;
wire            n1735____DOLLAR__4585;
wire            n1736____DOLLAR__4586;
wire            n1737____DOLLAR__4587;
wire            n1738____DOLLAR__4588;
wire            n1739____DOLLAR__4589;
wire            n173____DOLLAR__761;
wire            n1740____DOLLAR__4590;
wire            n1741____DOLLAR__4591;
wire            n1742____DOLLAR__4592;
wire            n1743____DOLLAR__4593;
wire            n1744____DOLLAR__4594;
wire            n1745____DOLLAR__4595;
wire            n1746____DOLLAR__4596;
wire            n1747____DOLLAR__4597;
wire            n1748____DOLLAR__4598;
wire            n1749____DOLLAR__4599;
wire            n174____DOLLAR__765;
wire            n1750____DOLLAR__4600;
wire            n1751____DOLLAR__4601;
wire            n1752____DOLLAR__4602;
wire            n1753____DOLLAR__4603;
wire            n1754____DOLLAR__4604;
wire            n1755____DOLLAR__4605;
wire            n1756____DOLLAR__4606;
wire            n1757____DOLLAR__4607;
wire            n1758____DOLLAR__4608;
wire            n1759____DOLLAR__4609;
wire            n175____DOLLAR__769;
wire            n1760____DOLLAR__4610;
wire            n1761____DOLLAR__4611;
wire            n1762____DOLLAR__4612;
wire            n1763____DOLLAR__4613;
wire            n1764____DOLLAR__4614;
wire            n1765____DOLLAR__4615;
wire            n1766____DOLLAR__4616;
wire            n1767____DOLLAR__4617;
wire            n1768____DOLLAR__4618;
wire            n1769____DOLLAR__4619;
wire            n176____DOLLAR__773;
wire            n1770____DOLLAR__4620;
wire            n1771____DOLLAR__4621;
wire            n1772____DOLLAR__4622;
wire            n1773____DOLLAR__4623;
wire            n1774____DOLLAR__4624;
wire            n1775____DOLLAR__4625;
wire            n1776____DOLLAR__4626;
wire            n1777____DOLLAR__4627;
wire            n1778____DOLLAR__4628;
wire            n1779____DOLLAR__4629;
wire            n177____DOLLAR__777;
wire            n1780____DOLLAR__4630;
wire            n1781____DOLLAR__4631;
wire            n1782____DOLLAR__4632;
wire            n1783____DOLLAR__4633;
wire            n1784____DOLLAR__4634;
wire            n1785____DOLLAR__4635;
wire            n1786____DOLLAR__4636;
wire            n1787____DOLLAR__4637;
wire            n1788____DOLLAR__4638;
wire            n1789____DOLLAR__4639;
wire            n178____DOLLAR__781;
wire            n1790____DOLLAR__4640;
wire            n1791____DOLLAR__4641;
wire            n1792____DOLLAR__4642;
wire            n1793____DOLLAR__4643;
wire            n1794____DOLLAR__4644;
wire            n1795____DOLLAR__4645;
wire            n1796____DOLLAR__4646;
wire            n1797____DOLLAR__4647;
wire            n1798____DOLLAR__4648;
wire            n1799____DOLLAR__4649;
wire            n179____DOLLAR__785;
wire            n17____DOLLAR__137;
wire            n1800____DOLLAR__4650;
wire            n1801____DOLLAR__4651;
wire            n1802____DOLLAR__4652;
wire            n1803____DOLLAR__4653;
wire            n1804____DOLLAR__4654;
wire            n1805____DOLLAR__4655;
wire            n1806____DOLLAR__4656;
wire            n1807____DOLLAR__4657;
wire            n1808____DOLLAR__4658;
wire            n1809____DOLLAR__4659;
wire            n180____DOLLAR__789;
wire            n1810____DOLLAR__4660;
wire            n1811____DOLLAR__4661;
wire            n1812____DOLLAR__4662;
wire            n1813____DOLLAR__4663;
wire            n1814____DOLLAR__4664;
wire            n1815____DOLLAR__4665;
wire            n1816____DOLLAR__4666;
wire            n1817____DOLLAR__4667;
wire            n1818____DOLLAR__4668;
wire            n1819____DOLLAR__4669;
wire            n181____DOLLAR__793;
wire            n1820____DOLLAR__4670;
wire            n1821____DOLLAR__4671;
wire            n1822____DOLLAR__4672;
wire            n1823____DOLLAR__4673;
wire            n1824____DOLLAR__4674;
wire            n1825____DOLLAR__4675;
wire            n1826____DOLLAR__4676;
wire            n1827____DOLLAR__4677;
wire            n1828____DOLLAR__4678;
wire            n1829____DOLLAR__4679;
wire            n182____DOLLAR__797;
wire            n1830____DOLLAR__4680;
wire            n1831____DOLLAR__4681;
wire            n1832____DOLLAR__4682;
wire            n1833____DOLLAR__4683;
wire            n1834____DOLLAR__4684;
wire            n1835____DOLLAR__4685;
wire            n1836____DOLLAR__4686;
wire            n1837____DOLLAR__4687;
wire            n1838____DOLLAR__4688;
wire            n1839____DOLLAR__4689;
wire            n183____DOLLAR__801;
wire            n1840____DOLLAR__4690;
wire            n1841____DOLLAR__4691;
wire            n1842____DOLLAR__4692;
wire            n1843____DOLLAR__4693;
wire            n1844____DOLLAR__4694;
wire            n1845____DOLLAR__4695;
wire            n1846____DOLLAR__4696;
wire            n1847____DOLLAR__4697;
wire            n1848____DOLLAR__4698;
wire            n1849____DOLLAR__4699;
wire            n184____DOLLAR__805;
wire            n1850____DOLLAR__4700;
wire            n1851____DOLLAR__4701;
wire            n1852____DOLLAR__4702;
wire            n1853____DOLLAR__4703;
wire            n1854____DOLLAR__4704;
wire            n1855____DOLLAR__4705;
wire            n1856____DOLLAR__4706;
wire            n1857____DOLLAR__4707;
wire            n1858____DOLLAR__4708;
wire            n1859____DOLLAR__4709;
wire            n185____DOLLAR__809;
wire            n1860____DOLLAR__4710;
wire            n1861____DOLLAR__4711;
wire            n1862____DOLLAR__4712;
wire            n1863____DOLLAR__4713;
wire            n1864____DOLLAR__4714;
wire            n1865____DOLLAR__4715;
wire            n1866____DOLLAR__4716;
wire            n1867____DOLLAR__4717;
wire            n1868____DOLLAR__4718;
wire            n1869____DOLLAR__4719;
wire            n186____DOLLAR__813;
wire            n1870____DOLLAR__4720;
wire            n1871____DOLLAR__4721;
wire            n1872____DOLLAR__4722;
wire            n1873____DOLLAR__4723;
wire            n1874____DOLLAR__4724;
wire            n1875____DOLLAR__4725;
wire            n1876____DOLLAR__4726;
wire            n1877____DOLLAR__4727;
wire            n1878____DOLLAR__4728;
wire            n1879____DOLLAR__4729;
wire            n187____DOLLAR__817;
wire            n1880____DOLLAR__4730;
wire            n1881____DOLLAR__4731;
wire            n1882____DOLLAR__4732;
wire            n1883____DOLLAR__4733;
wire            n1884____DOLLAR__4734;
wire            n1885____DOLLAR__4735;
wire            n1886____DOLLAR__4736;
wire            n1887____DOLLAR__4737;
wire            n1888____DOLLAR__4738;
wire            n1889____DOLLAR__4739;
wire            n188____DOLLAR__821;
wire            n1890____DOLLAR__4740;
wire            n1891____DOLLAR__4741;
wire            n1892____DOLLAR__4742;
wire            n1893____DOLLAR__4743;
wire            n1894____DOLLAR__4744;
wire            n1895____DOLLAR__4745;
wire            n1896____DOLLAR__4746;
wire            n1897____DOLLAR__4747;
wire            n1898____DOLLAR__4748;
wire            n1899____DOLLAR__4749;
wire            n189____DOLLAR__825;
wire            n18____DOLLAR__141;
wire            n1900____DOLLAR__4750;
wire            n1901____DOLLAR__4751;
wire            n1902____DOLLAR__4752;
wire            n1903____DOLLAR__4753;
wire            n1904____DOLLAR__4754;
wire            n1905____DOLLAR__4755;
wire            n1906____DOLLAR__4756;
wire            n1907____DOLLAR__4757;
wire            n1908____DOLLAR__4758;
wire            n1909____DOLLAR__4759;
wire            n190____DOLLAR__829;
wire            n1910____DOLLAR__4760;
wire            n1911____DOLLAR__4761;
wire            n1912____DOLLAR__4762;
wire            n1913____DOLLAR__4763;
wire            n1914____DOLLAR__4764;
wire            n1915____DOLLAR__4765;
wire            n1916____DOLLAR__4766;
wire            n1917____DOLLAR__4767;
wire            n1918____DOLLAR__4768;
wire            n1919____DOLLAR__4769;
wire            n191____DOLLAR__833;
wire            n1920____DOLLAR__4770;
wire            n1921____DOLLAR__4771;
wire            n1922____DOLLAR__4772;
wire            n1923____DOLLAR__4773;
wire            n1924____DOLLAR__4774;
wire            n1925____DOLLAR__4775;
wire            n1926____DOLLAR__4776;
wire            n1927____DOLLAR__4777;
wire            n1928____DOLLAR__4778;
wire            n1929____DOLLAR__4779;
wire            n192____DOLLAR__837;
wire            n1930____DOLLAR__4780;
wire            n1931____DOLLAR__4781;
wire            n1932____DOLLAR__4782;
wire            n1933____DOLLAR__4783;
wire            n1934____DOLLAR__4784;
wire            n1935____DOLLAR__4785;
wire            n1936____DOLLAR__4786;
wire            n1937____DOLLAR__4787;
wire            n1938____DOLLAR__4788;
wire            n1939____DOLLAR__4789;
wire            n193____DOLLAR__841;
wire            n1940____DOLLAR__4790;
wire            n1941____DOLLAR__4791;
wire            n1942____DOLLAR__4792;
wire            n1943____DOLLAR__4793;
wire            n1944____DOLLAR__4794;
wire            n1945____DOLLAR__4795;
wire            n1946____DOLLAR__4796;
wire            n1947____DOLLAR__4797;
wire            n1948____DOLLAR__4798;
wire            n1949____DOLLAR__4799;
wire            n194____DOLLAR__845;
wire            n1950____DOLLAR__4800;
wire            n1951____DOLLAR__4801;
wire            n1952____DOLLAR__4802;
wire            n1953____DOLLAR__4808;
wire            n1954____DOLLAR__4812;
wire      [4:0] n1955____DOLLAR__4814;
wire      [7:0] n1956____DOLLAR__4822;
wire      [7:0] n1957____DOLLAR__4824;
wire      [7:0] n1958____DOLLAR__4828;
wire      [7:0] n1959____DOLLAR__4829;
wire            n195____DOLLAR__849;
wire            n1960____DOLLAR__4832;
wire      [2:0] n1961____DOLLAR__4839;
wire      [7:0] n1962____DOLLAR__4841;
wire      [7:0] n1963____DOLLAR__4843;
wire      [7:0] n1964____DOLLAR__4844;
wire            n1965____DOLLAR__4848;
wire            n1966____DOLLAR__4850;
wire      [4:0] n1967____DOLLAR__4852;
wire      [7:0] n1968____DOLLAR__4858;
wire      [7:0] n1969____DOLLAR__4860;
wire            n196____DOLLAR__853;
wire      [7:0] n1970____DOLLAR__4862;
wire      [7:0] n1971____DOLLAR__4863;
wire            n1972____DOLLAR__4864;
wire            n1973____DOLLAR__4868;
wire            n1974____DOLLAR__4873;
wire            n1975____DOLLAR__4875;
wire      [4:0] n1976____DOLLAR__4880;
wire      [7:0] n1977____DOLLAR__4886;
wire      [4:0] n1978____DOLLAR__4891;
wire      [7:0] n1979____DOLLAR__4893;
wire            n197____DOLLAR__857;
wire      [7:0] n1980____DOLLAR__4895;
wire      [7:0] n1981____DOLLAR__4896;
wire      [3:0] n1982____DOLLAR__187085;
wire            n1983____DOLLAR__187166;
wire            n1984____DOLLAR__187161;
wire            n1985____DOLLAR__187156;
wire            n1986____DOLLAR__187151;
wire            n1987____DOLLAR__187146;
wire            n1988____DOLLAR__187141;
wire            n1989____DOLLAR__187136;
wire            n198____DOLLAR__861;
wire            n1990____DOLLAR__187131;
wire            n1991____DOLLAR__187126;
wire            n1992____DOLLAR__187121;
wire            n1993____DOLLAR__187116;
wire            n1994____DOLLAR__187111;
wire            n1995____DOLLAR__187106;
wire            n1996____DOLLAR__187101;
wire            n1997____DOLLAR__187096;
wire            n1998____DOLLAR__187091;
wire      [7:0] n1999____DOLLAR__187093;
wire            n199____DOLLAR__865;
wire            n19____DOLLAR__145;
wire      [7:0] n2000____DOLLAR__187098;
wire      [7:0] n2001____DOLLAR__187103;
wire      [7:0] n2002____DOLLAR__187108;
wire      [7:0] n2003____DOLLAR__187113;
wire      [7:0] n2004____DOLLAR__187118;
wire      [7:0] n2005____DOLLAR__187123;
wire      [7:0] n2006____DOLLAR__187128;
wire      [7:0] n2007____DOLLAR__187133;
wire      [7:0] n2008____DOLLAR__187138;
wire      [7:0] n2009____DOLLAR__187143;
wire            n200____DOLLAR__869;
wire      [7:0] n2010____DOLLAR__187148;
wire      [7:0] n2011____DOLLAR__187153;
wire      [7:0] n2012____DOLLAR__187158;
wire      [7:0] n2013____DOLLAR__187163;
wire      [7:0] n2014____DOLLAR__187168;
wire            n2015____DOLLAR__4902;
wire            n2016____DOLLAR__4904;
wire      [4:0] n2017____DOLLAR__4906;
wire      [7:0] n2018____DOLLAR__4912;
wire      [7:0] n2019____DOLLAR__4914;
wire            n201____DOLLAR__873;
wire      [7:0] n2020____DOLLAR__4916;
wire      [7:0] n2021____DOLLAR__4917;
wire            n2022____DOLLAR__4920;
wire            n2023____DOLLAR__4925;
wire            n2024____DOLLAR__4927;
wire      [4:0] n2025____DOLLAR__4929;
wire      [7:0] n2026____DOLLAR__4935;
wire      [7:0] n2027____DOLLAR__4937;
wire      [7:0] n2028____DOLLAR__4939;
wire      [7:0] n2029____DOLLAR__4940;
wire            n202____DOLLAR__877;
wire            n2030____DOLLAR__4943;
wire            n2031____DOLLAR__4948;
wire            n2032____DOLLAR__4950;
wire      [4:0] n2033____DOLLAR__4952;
wire      [7:0] n2034____DOLLAR__4958;
wire      [7:0] n2035____DOLLAR__4960;
wire      [7:0] n2036____DOLLAR__4962;
wire      [7:0] n2037____DOLLAR__4963;
wire            n2038____DOLLAR__4966;
wire            n2039____DOLLAR__4971;
wire            n203____DOLLAR__881;
wire            n2040____DOLLAR__4973;
wire      [4:0] n2041____DOLLAR__4975;
wire      [7:0] n2042____DOLLAR__4981;
wire      [7:0] n2043____DOLLAR__4983;
wire      [7:0] n2044____DOLLAR__4985;
wire      [7:0] n2045____DOLLAR__4986;
wire            n2046____DOLLAR__4989;
wire            n2047____DOLLAR__4994;
wire            n2048____DOLLAR__4996;
wire      [4:0] n2049____DOLLAR__4998;
wire            n204____DOLLAR__885;
wire      [7:0] n2050____DOLLAR__5004;
wire      [7:0] n2051____DOLLAR__5006;
wire      [7:0] n2052____DOLLAR__5008;
wire      [7:0] n2053____DOLLAR__5009;
wire            n2054____DOLLAR__5012;
wire            n2055____DOLLAR__5017;
wire            n2056____DOLLAR__5019;
wire      [4:0] n2057____DOLLAR__5021;
wire      [7:0] n2058____DOLLAR__5027;
wire      [7:0] n2059____DOLLAR__5029;
wire            n205____DOLLAR__889;
wire      [7:0] n2060____DOLLAR__5031;
wire      [7:0] n2061____DOLLAR__5032;
wire            n2062____DOLLAR__5035;
wire            n2063____DOLLAR__5040;
wire            n2064____DOLLAR__5042;
wire      [4:0] n2065____DOLLAR__5044;
wire      [7:0] n2066____DOLLAR__5050;
wire      [7:0] n2067____DOLLAR__5052;
wire      [7:0] n2068____DOLLAR__5054;
wire      [7:0] n2069____DOLLAR__5055;
wire            n206____DOLLAR__893;
wire            n2070____DOLLAR__5058;
wire            n2071____DOLLAR__5063;
wire            n2072____DOLLAR__5065;
wire      [4:0] n2073____DOLLAR__5067;
wire      [7:0] n2074____DOLLAR__5073;
wire      [7:0] n2075____DOLLAR__5075;
wire      [7:0] n2076____DOLLAR__5077;
wire      [7:0] n2077____DOLLAR__5078;
wire            n2078____DOLLAR__5081;
wire            n2079____DOLLAR__5086;
wire            n207____DOLLAR__897;
wire            n2080____DOLLAR__5088;
wire      [4:0] n2081____DOLLAR__5090;
wire      [7:0] n2082____DOLLAR__5096;
wire      [7:0] n2083____DOLLAR__5098;
wire      [7:0] n2084____DOLLAR__5100;
wire      [7:0] n2085____DOLLAR__5101;
wire            n2086____DOLLAR__5104;
wire            n2087____DOLLAR__5109;
wire            n2088____DOLLAR__5111;
wire      [4:0] n2089____DOLLAR__5113;
wire            n208____DOLLAR__901;
wire      [7:0] n2090____DOLLAR__5119;
wire      [7:0] n2091____DOLLAR__5121;
wire      [7:0] n2092____DOLLAR__5123;
wire      [7:0] n2093____DOLLAR__5124;
wire            n2094____DOLLAR__5127;
wire            n2095____DOLLAR__5132;
wire            n2096____DOLLAR__5134;
wire      [4:0] n2097____DOLLAR__5136;
wire      [7:0] n2098____DOLLAR__5142;
wire      [7:0] n2099____DOLLAR__5144;
wire            n209____DOLLAR__905;
wire            n20____DOLLAR__149;
wire      [7:0] n2100____DOLLAR__5146;
wire      [7:0] n2101____DOLLAR__5147;
wire            n2102____DOLLAR__5150;
wire            n2103____DOLLAR__5155;
wire            n2104____DOLLAR__5157;
wire      [4:0] n2105____DOLLAR__5159;
wire      [7:0] n2106____DOLLAR__5165;
wire      [7:0] n2107____DOLLAR__5167;
wire      [7:0] n2108____DOLLAR__5169;
wire      [7:0] n2109____DOLLAR__5170;
wire            n210____DOLLAR__909;
wire            n2110____DOLLAR__5173;
wire            n2111____DOLLAR__5178;
wire            n2112____DOLLAR__5180;
wire      [4:0] n2113____DOLLAR__5182;
wire      [7:0] n2114____DOLLAR__5188;
wire      [7:0] n2115____DOLLAR__5190;
wire      [7:0] n2116____DOLLAR__5192;
wire      [7:0] n2117____DOLLAR__5193;
wire            n2118____DOLLAR__5196;
wire            n2119____DOLLAR__5201;
wire            n211____DOLLAR__913;
wire            n2120____DOLLAR__5203;
wire      [4:0] n2121____DOLLAR__5205;
wire      [7:0] n2122____DOLLAR__5211;
wire      [7:0] n2123____DOLLAR__5213;
wire      [7:0] n2124____DOLLAR__5215;
wire      [7:0] n2125____DOLLAR__5216;
wire            n2126____DOLLAR__5219;
wire            n2127____DOLLAR__5224;
wire            n2128____DOLLAR__5226;
wire      [4:0] n2129____DOLLAR__5228;
wire            n212____DOLLAR__917;
wire      [7:0] n2130____DOLLAR__5234;
wire      [7:0] n2131____DOLLAR__5236;
wire      [7:0] n2132____DOLLAR__5238;
wire      [7:0] n2133____DOLLAR__5239;
wire            n2134____DOLLAR__5242;
wire            n2135____DOLLAR__5247;
wire            n2136____DOLLAR__5249;
wire      [4:0] n2137____DOLLAR__5251;
wire      [7:0] n2138____DOLLAR__5257;
wire      [7:0] n2139____DOLLAR__5259;
wire            n213____DOLLAR__921;
wire      [7:0] n2140____DOLLAR__5261;
wire      [7:0] n2141____DOLLAR__5262;
wire            n2142____DOLLAR__5265;
wire            n2143____DOLLAR__5270;
wire            n2144____DOLLAR__5272;
wire      [4:0] n2145____DOLLAR__5274;
wire      [7:0] n2146____DOLLAR__5280;
wire      [7:0] n2147____DOLLAR__5282;
wire      [7:0] n2148____DOLLAR__5284;
wire      [7:0] n2149____DOLLAR__5285;
wire            n214____DOLLAR__925;
wire            n2150____DOLLAR__5288;
wire            n2151____DOLLAR__5293;
wire            n2152____DOLLAR__5295;
wire      [4:0] n2153____DOLLAR__5297;
wire      [7:0] n2154____DOLLAR__5303;
wire      [7:0] n2155____DOLLAR__5305;
wire      [7:0] n2156____DOLLAR__5307;
wire      [7:0] n2157____DOLLAR__5308;
wire            n2158____DOLLAR__5311;
wire            n2159____DOLLAR__5316;
wire            n215____DOLLAR__929;
wire            n2160____DOLLAR__5318;
wire      [4:0] n2161____DOLLAR__5320;
wire      [7:0] n2162____DOLLAR__5326;
wire      [7:0] n2163____DOLLAR__5328;
wire      [7:0] n2164____DOLLAR__5330;
wire      [7:0] n2165____DOLLAR__5331;
wire            n2166____DOLLAR__5334;
wire            n2167____DOLLAR__5339;
wire            n2168____DOLLAR__5341;
wire      [4:0] n2169____DOLLAR__5343;
wire            n216____DOLLAR__933;
wire      [7:0] n2170____DOLLAR__5349;
wire      [7:0] n2171____DOLLAR__5351;
wire      [7:0] n2172____DOLLAR__5353;
wire      [7:0] n2173____DOLLAR__5354;
wire            n2174____DOLLAR__5357;
wire            n2175____DOLLAR__5362;
wire            n2176____DOLLAR__5364;
wire      [4:0] n2177____DOLLAR__5366;
wire      [7:0] n2178____DOLLAR__5372;
wire      [7:0] n2179____DOLLAR__5374;
wire            n217____DOLLAR__937;
wire      [7:0] n2180____DOLLAR__5376;
wire      [7:0] n2181____DOLLAR__5377;
wire            n2182____DOLLAR__5380;
wire      [7:0] n2183____DOLLAR__5384;
wire      [7:0] n2184____DOLLAR__5385;
wire      [7:0] n2185____DOLLAR__5386;
wire      [7:0] n2186____DOLLAR__5387;
wire      [7:0] n2187____DOLLAR__5388;
wire      [7:0] n2188____DOLLAR__5389;
wire      [7:0] n2189____DOLLAR__5390;
wire            n218____DOLLAR__941;
wire      [7:0] n2190____DOLLAR__5391;
wire      [7:0] n2191____DOLLAR__5392;
wire      [7:0] n2192____DOLLAR__5393;
wire      [7:0] n2193____DOLLAR__5394;
wire      [7:0] n2194____DOLLAR__5395;
wire      [7:0] n2195____DOLLAR__5396;
wire      [7:0] n2196____DOLLAR__5397;
wire      [7:0] n2197____DOLLAR__5398;
wire      [7:0] n2198____DOLLAR__5399;
wire      [7:0] n2199____DOLLAR__5400;
wire            n219____DOLLAR__945;
wire            n21____DOLLAR__153;
wire      [7:0] n2200____DOLLAR__5401;
wire      [7:0] n2201____DOLLAR__5402;
wire      [7:0] n2202____DOLLAR__5403;
wire      [7:0] n2203____DOLLAR__5404;
wire      [7:0] n2204____DOLLAR__5405;
wire      [7:0] n2205____DOLLAR__5406;
wire            n2206____DOLLAR__5407;
wire      [7:0] n2207____DOLLAR__5409;
wire      [2:0] n2208____DOLLAR__5414;
wire      [7:0] n2209____DOLLAR__5416;
wire            n220____DOLLAR__949;
wire      [7:0] n2210____DOLLAR__5418;
wire      [7:0] n2211____DOLLAR__5419;
wire      [7:0] n2212____DOLLAR__5420;
wire      [7:0] n2213____DOLLAR__5421;
wire            n2214____DOLLAR__5426;
wire            n2215____DOLLAR__5430;
wire            n2216____DOLLAR__5432;
wire      [1:0] n2217____DOLLAR__5437;
wire      [4:0] n2218____DOLLAR__5445;
wire      [7:0] n2219____DOLLAR__5451;
wire            n221____DOLLAR__953;
wire      [3:0] n2220____DOLLAR__192041;
wire            n2221____DOLLAR__192122;
wire            n2222____DOLLAR__192117;
wire            n2223____DOLLAR__192112;
wire            n2224____DOLLAR__192107;
wire            n2225____DOLLAR__192102;
wire            n2226____DOLLAR__192097;
wire            n2227____DOLLAR__192092;
wire            n2228____DOLLAR__192087;
wire            n2229____DOLLAR__192082;
wire            n222____DOLLAR__957;
wire            n2230____DOLLAR__192077;
wire            n2231____DOLLAR__192072;
wire            n2232____DOLLAR__192067;
wire            n2233____DOLLAR__192062;
wire            n2234____DOLLAR__192057;
wire            n2235____DOLLAR__192052;
wire            n2236____DOLLAR__192047;
wire      [7:0] n2237____DOLLAR__192049;
wire      [7:0] n2238____DOLLAR__192054;
wire      [7:0] n2239____DOLLAR__192059;
wire            n223____DOLLAR__961;
wire      [7:0] n2240____DOLLAR__192064;
wire      [7:0] n2241____DOLLAR__192069;
wire      [7:0] n2242____DOLLAR__192074;
wire      [7:0] n2243____DOLLAR__192079;
wire      [7:0] n2244____DOLLAR__192084;
wire      [7:0] n2245____DOLLAR__192089;
wire      [7:0] n2246____DOLLAR__192094;
wire      [7:0] n2247____DOLLAR__192099;
wire      [7:0] n2248____DOLLAR__192104;
wire      [7:0] n2249____DOLLAR__192109;
wire            n224____DOLLAR__965;
wire      [7:0] n2250____DOLLAR__192114;
wire      [7:0] n2251____DOLLAR__192119;
wire      [7:0] n2252____DOLLAR__192124;
wire     [15:0] n2253____DOLLAR__5459;
wire            n2254____DOLLAR__5465;
wire            n2255____DOLLAR__5469;
wire            n2256____DOLLAR__5471;
wire      [1:0] n2257____DOLLAR__5476;
wire      [4:0] n2258____DOLLAR__5484;
wire      [7:0] n2259____DOLLAR__5490;
wire            n225____DOLLAR__969;
wire      [3:0] n2260____DOLLAR__192149;
wire            n2261____DOLLAR__192230;
wire            n2262____DOLLAR__192225;
wire            n2263____DOLLAR__192220;
wire            n2264____DOLLAR__192215;
wire            n2265____DOLLAR__192210;
wire            n2266____DOLLAR__192205;
wire            n2267____DOLLAR__192200;
wire            n2268____DOLLAR__192195;
wire            n2269____DOLLAR__192190;
wire            n226____DOLLAR__973;
wire            n2270____DOLLAR__192185;
wire            n2271____DOLLAR__192180;
wire            n2272____DOLLAR__192175;
wire            n2273____DOLLAR__192170;
wire            n2274____DOLLAR__192165;
wire            n2275____DOLLAR__192160;
wire            n2276____DOLLAR__192155;
wire      [7:0] n2277____DOLLAR__192157;
wire      [7:0] n2278____DOLLAR__192162;
wire      [7:0] n2279____DOLLAR__192167;
wire            n227____DOLLAR__977;
wire      [7:0] n2280____DOLLAR__192172;
wire      [7:0] n2281____DOLLAR__192177;
wire      [7:0] n2282____DOLLAR__192182;
wire      [7:0] n2283____DOLLAR__192187;
wire      [7:0] n2284____DOLLAR__192192;
wire      [7:0] n2285____DOLLAR__192197;
wire      [7:0] n2286____DOLLAR__192202;
wire      [7:0] n2287____DOLLAR__192207;
wire      [7:0] n2288____DOLLAR__192212;
wire      [7:0] n2289____DOLLAR__192217;
wire            n228____DOLLAR__981;
wire      [7:0] n2290____DOLLAR__192222;
wire      [7:0] n2291____DOLLAR__192227;
wire      [7:0] n2292____DOLLAR__192232;
wire     [15:0] n2293____DOLLAR__5498;
wire            n2294____DOLLAR__5504;
wire            n2295____DOLLAR__5508;
wire            n2296____DOLLAR__5510;
wire     [15:0] n2297____DOLLAR__5515;
wire            n2298____DOLLAR__5521;
wire            n2299____DOLLAR__5525;
wire            n229____DOLLAR__985;
wire            n22____DOLLAR__157;
wire            n2300____DOLLAR__5529;
wire            n2301____DOLLAR__5533;
wire            n2302____DOLLAR__5537;
wire            n2303____DOLLAR__5541;
wire            n2304____DOLLAR__5545;
wire            n2305____DOLLAR__5549;
wire            n2306____DOLLAR__5553;
wire            n2307____DOLLAR__5557;
wire            n2308____DOLLAR__5561;
wire            n2309____DOLLAR__5565;
wire            n230____DOLLAR__989;
wire            n2310____DOLLAR__5569;
wire            n2311____DOLLAR__5573;
wire            n2312____DOLLAR__5577;
wire            n2313____DOLLAR__5581;
wire            n2314____DOLLAR__5585;
wire            n2315____DOLLAR__5589;
wire            n2316____DOLLAR__5593;
wire            n2317____DOLLAR__5597;
wire            n2318____DOLLAR__5601;
wire            n2319____DOLLAR__5605;
wire            n231____DOLLAR__993;
wire            n2320____DOLLAR__5609;
wire            n2321____DOLLAR__5613;
wire            n2322____DOLLAR__5617;
wire            n2323____DOLLAR__5621;
wire            n2324____DOLLAR__5625;
wire            n2325____DOLLAR__5629;
wire            n2326____DOLLAR__5633;
wire            n2327____DOLLAR__5637;
wire            n2328____DOLLAR__5641;
wire            n2329____DOLLAR__5645;
wire            n232____DOLLAR__995;
wire            n2330____DOLLAR__5649;
wire            n2331____DOLLAR__5653;
wire            n2332____DOLLAR__5657;
wire            n2333____DOLLAR__5661;
wire            n2334____DOLLAR__5665;
wire            n2335____DOLLAR__5669;
wire            n2336____DOLLAR__5673;
wire            n2337____DOLLAR__5677;
wire            n2338____DOLLAR__5681;
wire            n2339____DOLLAR__5685;
wire            n233____DOLLAR__996;
wire            n2340____DOLLAR__5689;
wire            n2341____DOLLAR__5693;
wire            n2342____DOLLAR__5697;
wire            n2343____DOLLAR__5701;
wire            n2344____DOLLAR__5705;
wire            n2345____DOLLAR__5709;
wire            n2346____DOLLAR__5713;
wire            n2347____DOLLAR__5717;
wire            n2348____DOLLAR__5721;
wire            n2349____DOLLAR__5725;
wire            n234____DOLLAR__997;
wire            n2350____DOLLAR__5729;
wire            n2351____DOLLAR__5733;
wire            n2352____DOLLAR__5737;
wire            n2353____DOLLAR__5741;
wire            n2354____DOLLAR__5745;
wire            n2355____DOLLAR__5749;
wire            n2356____DOLLAR__5753;
wire            n2357____DOLLAR__5757;
wire            n2358____DOLLAR__5761;
wire            n2359____DOLLAR__5765;
wire            n235____DOLLAR__998;
wire            n2360____DOLLAR__5769;
wire            n2361____DOLLAR__5773;
wire            n2362____DOLLAR__5777;
wire            n2363____DOLLAR__5781;
wire            n2364____DOLLAR__5785;
wire            n2365____DOLLAR__5789;
wire            n2366____DOLLAR__5793;
wire            n2367____DOLLAR__5797;
wire            n2368____DOLLAR__5801;
wire            n2369____DOLLAR__5805;
wire            n236____DOLLAR__999;
wire            n2370____DOLLAR__5809;
wire            n2371____DOLLAR__5813;
wire            n2372____DOLLAR__5817;
wire            n2373____DOLLAR__5821;
wire            n2374____DOLLAR__5825;
wire            n2375____DOLLAR__5829;
wire            n2376____DOLLAR__5833;
wire            n2377____DOLLAR__5837;
wire            n2378____DOLLAR__5841;
wire            n2379____DOLLAR__5845;
wire            n237____DOLLAR__1000;
wire            n2380____DOLLAR__5849;
wire            n2381____DOLLAR__5853;
wire            n2382____DOLLAR__5857;
wire            n2383____DOLLAR__5861;
wire            n2384____DOLLAR__5865;
wire            n2385____DOLLAR__5869;
wire            n2386____DOLLAR__5873;
wire            n2387____DOLLAR__5877;
wire            n2388____DOLLAR__5881;
wire            n2389____DOLLAR__5885;
wire            n238____DOLLAR__1001;
wire            n2390____DOLLAR__5889;
wire            n2391____DOLLAR__5893;
wire            n2392____DOLLAR__5897;
wire            n2393____DOLLAR__5901;
wire            n2394____DOLLAR__5905;
wire            n2395____DOLLAR__5909;
wire            n2396____DOLLAR__5913;
wire            n2397____DOLLAR__5917;
wire            n2398____DOLLAR__5921;
wire            n2399____DOLLAR__5925;
wire            n239____DOLLAR__1002;
wire            n23____DOLLAR__161;
wire            n2400____DOLLAR__5929;
wire            n2401____DOLLAR__5933;
wire            n2402____DOLLAR__5937;
wire            n2403____DOLLAR__5941;
wire            n2404____DOLLAR__5945;
wire            n2405____DOLLAR__5949;
wire            n2406____DOLLAR__5953;
wire            n2407____DOLLAR__5957;
wire            n2408____DOLLAR__5961;
wire            n2409____DOLLAR__5965;
wire            n240____DOLLAR__1003;
wire            n2410____DOLLAR__5969;
wire            n2411____DOLLAR__5973;
wire            n2412____DOLLAR__5977;
wire            n2413____DOLLAR__5981;
wire            n2414____DOLLAR__5985;
wire            n2415____DOLLAR__5989;
wire            n2416____DOLLAR__5993;
wire            n2417____DOLLAR__5997;
wire            n2418____DOLLAR__6001;
wire            n2419____DOLLAR__6005;
wire            n241____DOLLAR__1004;
wire            n2420____DOLLAR__6009;
wire            n2421____DOLLAR__6013;
wire            n2422____DOLLAR__6017;
wire            n2423____DOLLAR__6021;
wire            n2424____DOLLAR__6025;
wire            n2425____DOLLAR__6029;
wire            n2426____DOLLAR__6033;
wire            n2427____DOLLAR__6037;
wire            n2428____DOLLAR__6041;
wire            n2429____DOLLAR__6045;
wire            n242____DOLLAR__1005;
wire            n2430____DOLLAR__6049;
wire            n2431____DOLLAR__6053;
wire            n2432____DOLLAR__6057;
wire            n2433____DOLLAR__6061;
wire            n2434____DOLLAR__6065;
wire            n2435____DOLLAR__6069;
wire            n2436____DOLLAR__6073;
wire            n2437____DOLLAR__6077;
wire            n2438____DOLLAR__6081;
wire            n2439____DOLLAR__6085;
wire            n243____DOLLAR__1006;
wire            n2440____DOLLAR__6089;
wire            n2441____DOLLAR__6093;
wire            n2442____DOLLAR__6097;
wire            n2443____DOLLAR__6101;
wire            n2444____DOLLAR__6105;
wire            n2445____DOLLAR__6109;
wire            n2446____DOLLAR__6113;
wire            n2447____DOLLAR__6117;
wire            n2448____DOLLAR__6121;
wire            n2449____DOLLAR__6125;
wire            n244____DOLLAR__1007;
wire            n2450____DOLLAR__6129;
wire            n2451____DOLLAR__6133;
wire            n2452____DOLLAR__6137;
wire            n2453____DOLLAR__6141;
wire            n2454____DOLLAR__6145;
wire            n2455____DOLLAR__6149;
wire            n2456____DOLLAR__6153;
wire            n2457____DOLLAR__6157;
wire            n2458____DOLLAR__6161;
wire            n2459____DOLLAR__6165;
wire            n245____DOLLAR__1008;
wire            n2460____DOLLAR__6169;
wire            n2461____DOLLAR__6173;
wire            n2462____DOLLAR__6177;
wire            n2463____DOLLAR__6181;
wire            n2464____DOLLAR__6185;
wire            n2465____DOLLAR__6189;
wire            n2466____DOLLAR__6193;
wire            n2467____DOLLAR__6197;
wire            n2468____DOLLAR__6201;
wire            n2469____DOLLAR__6205;
wire            n246____DOLLAR__1009;
wire            n2470____DOLLAR__6209;
wire            n2471____DOLLAR__6213;
wire            n2472____DOLLAR__6217;
wire            n2473____DOLLAR__6221;
wire            n2474____DOLLAR__6225;
wire            n2475____DOLLAR__6229;
wire            n2476____DOLLAR__6233;
wire            n2477____DOLLAR__6237;
wire            n2478____DOLLAR__6241;
wire            n2479____DOLLAR__6245;
wire            n247____DOLLAR__1010;
wire            n2480____DOLLAR__6249;
wire            n2481____DOLLAR__6253;
wire            n2482____DOLLAR__6257;
wire            n2483____DOLLAR__6261;
wire            n2484____DOLLAR__6265;
wire            n2485____DOLLAR__6269;
wire            n2486____DOLLAR__6273;
wire            n2487____DOLLAR__6277;
wire            n2488____DOLLAR__6281;
wire            n2489____DOLLAR__6285;
wire            n248____DOLLAR__1011;
wire            n2490____DOLLAR__6289;
wire            n2491____DOLLAR__6293;
wire            n2492____DOLLAR__6297;
wire            n2493____DOLLAR__6301;
wire            n2494____DOLLAR__6305;
wire            n2495____DOLLAR__6309;
wire            n2496____DOLLAR__6313;
wire            n2497____DOLLAR__6317;
wire            n2498____DOLLAR__6321;
wire            n2499____DOLLAR__6325;
wire            n249____DOLLAR__1012;
wire            n24____DOLLAR__165;
wire            n2500____DOLLAR__6329;
wire            n2501____DOLLAR__6333;
wire            n2502____DOLLAR__6337;
wire            n2503____DOLLAR__6341;
wire            n2504____DOLLAR__6345;
wire            n2505____DOLLAR__6349;
wire            n2506____DOLLAR__6353;
wire            n2507____DOLLAR__6357;
wire            n2508____DOLLAR__6361;
wire            n2509____DOLLAR__6365;
wire            n250____DOLLAR__1013;
wire            n2510____DOLLAR__6369;
wire            n2511____DOLLAR__6373;
wire            n2512____DOLLAR__6377;
wire            n2513____DOLLAR__6381;
wire            n2514____DOLLAR__6385;
wire            n2515____DOLLAR__6389;
wire            n2516____DOLLAR__6393;
wire            n2517____DOLLAR__6397;
wire            n2518____DOLLAR__6401;
wire            n2519____DOLLAR__6405;
wire            n251____DOLLAR__1014;
wire            n2520____DOLLAR__6409;
wire            n2521____DOLLAR__6413;
wire            n2522____DOLLAR__6417;
wire            n2523____DOLLAR__6421;
wire            n2524____DOLLAR__6425;
wire            n2525____DOLLAR__6429;
wire            n2526____DOLLAR__6433;
wire            n2527____DOLLAR__6437;
wire            n2528____DOLLAR__6441;
wire            n2529____DOLLAR__6445;
wire            n252____DOLLAR__1015;
wire            n2530____DOLLAR__6449;
wire            n2531____DOLLAR__6453;
wire            n2532____DOLLAR__6457;
wire            n2533____DOLLAR__6461;
wire            n2534____DOLLAR__6465;
wire            n2535____DOLLAR__6469;
wire            n2536____DOLLAR__6473;
wire            n2537____DOLLAR__6477;
wire            n2538____DOLLAR__6481;
wire            n2539____DOLLAR__6485;
wire            n253____DOLLAR__1016;
wire            n2540____DOLLAR__6489;
wire            n2541____DOLLAR__6493;
wire            n2542____DOLLAR__6497;
wire            n2543____DOLLAR__6501;
wire            n2544____DOLLAR__6505;
wire            n2545____DOLLAR__6509;
wire            n2546____DOLLAR__6513;
wire            n2547____DOLLAR__6517;
wire            n2548____DOLLAR__6519;
wire            n2549____DOLLAR__6520;
wire            n254____DOLLAR__1017;
wire            n2550____DOLLAR__6521;
wire            n2551____DOLLAR__6522;
wire            n2552____DOLLAR__6523;
wire            n2553____DOLLAR__6524;
wire            n2554____DOLLAR__6525;
wire            n2555____DOLLAR__6526;
wire            n2556____DOLLAR__6527;
wire            n2557____DOLLAR__6528;
wire            n2558____DOLLAR__6529;
wire            n2559____DOLLAR__6530;
wire            n255____DOLLAR__1018;
wire            n2560____DOLLAR__6531;
wire            n2561____DOLLAR__6532;
wire            n2562____DOLLAR__6533;
wire            n2563____DOLLAR__6534;
wire            n2564____DOLLAR__6535;
wire            n2565____DOLLAR__6536;
wire            n2566____DOLLAR__6537;
wire            n2567____DOLLAR__6538;
wire            n2568____DOLLAR__6539;
wire            n2569____DOLLAR__6540;
wire            n256____DOLLAR__1019;
wire            n2570____DOLLAR__6541;
wire            n2571____DOLLAR__6542;
wire            n2572____DOLLAR__6543;
wire            n2573____DOLLAR__6544;
wire            n2574____DOLLAR__6545;
wire            n2575____DOLLAR__6546;
wire            n2576____DOLLAR__6547;
wire            n2577____DOLLAR__6548;
wire            n2578____DOLLAR__6549;
wire            n2579____DOLLAR__6550;
wire            n257____DOLLAR__1020;
wire            n2580____DOLLAR__6551;
wire            n2581____DOLLAR__6552;
wire            n2582____DOLLAR__6553;
wire            n2583____DOLLAR__6554;
wire            n2584____DOLLAR__6555;
wire            n2585____DOLLAR__6556;
wire            n2586____DOLLAR__6557;
wire            n2587____DOLLAR__6558;
wire            n2588____DOLLAR__6559;
wire            n2589____DOLLAR__6560;
wire            n258____DOLLAR__1021;
wire            n2590____DOLLAR__6561;
wire            n2591____DOLLAR__6562;
wire            n2592____DOLLAR__6563;
wire            n2593____DOLLAR__6564;
wire            n2594____DOLLAR__6565;
wire            n2595____DOLLAR__6566;
wire            n2596____DOLLAR__6567;
wire            n2597____DOLLAR__6568;
wire            n2598____DOLLAR__6569;
wire            n2599____DOLLAR__6570;
wire            n259____DOLLAR__1022;
wire            n25____DOLLAR__169;
wire            n2600____DOLLAR__6571;
wire            n2601____DOLLAR__6572;
wire            n2602____DOLLAR__6573;
wire            n2603____DOLLAR__6574;
wire            n2604____DOLLAR__6575;
wire            n2605____DOLLAR__6576;
wire            n2606____DOLLAR__6577;
wire            n2607____DOLLAR__6578;
wire            n2608____DOLLAR__6579;
wire            n2609____DOLLAR__6580;
wire            n260____DOLLAR__1023;
wire            n2610____DOLLAR__6581;
wire            n2611____DOLLAR__6582;
wire            n2612____DOLLAR__6583;
wire            n2613____DOLLAR__6584;
wire            n2614____DOLLAR__6585;
wire            n2615____DOLLAR__6586;
wire            n2616____DOLLAR__6587;
wire            n2617____DOLLAR__6588;
wire            n2618____DOLLAR__6589;
wire            n2619____DOLLAR__6590;
wire            n261____DOLLAR__1024;
wire            n2620____DOLLAR__6591;
wire            n2621____DOLLAR__6592;
wire            n2622____DOLLAR__6593;
wire            n2623____DOLLAR__6594;
wire            n2624____DOLLAR__6595;
wire            n2625____DOLLAR__6596;
wire            n2626____DOLLAR__6597;
wire            n2627____DOLLAR__6598;
wire            n2628____DOLLAR__6599;
wire            n2629____DOLLAR__6600;
wire            n262____DOLLAR__1025;
wire            n2630____DOLLAR__6601;
wire            n2631____DOLLAR__6602;
wire            n2632____DOLLAR__6603;
wire            n2633____DOLLAR__6604;
wire            n2634____DOLLAR__6605;
wire            n2635____DOLLAR__6606;
wire            n2636____DOLLAR__6607;
wire            n2637____DOLLAR__6608;
wire            n2638____DOLLAR__6609;
wire            n2639____DOLLAR__6610;
wire            n263____DOLLAR__1026;
wire            n2640____DOLLAR__6611;
wire            n2641____DOLLAR__6612;
wire            n2642____DOLLAR__6613;
wire            n2643____DOLLAR__6614;
wire            n2644____DOLLAR__6615;
wire            n2645____DOLLAR__6616;
wire            n2646____DOLLAR__6617;
wire            n2647____DOLLAR__6618;
wire            n2648____DOLLAR__6619;
wire            n2649____DOLLAR__6620;
wire            n264____DOLLAR__1027;
wire            n2650____DOLLAR__6621;
wire            n2651____DOLLAR__6622;
wire            n2652____DOLLAR__6623;
wire            n2653____DOLLAR__6624;
wire            n2654____DOLLAR__6625;
wire            n2655____DOLLAR__6626;
wire            n2656____DOLLAR__6627;
wire            n2657____DOLLAR__6628;
wire            n2658____DOLLAR__6629;
wire            n2659____DOLLAR__6630;
wire            n265____DOLLAR__1028;
wire            n2660____DOLLAR__6631;
wire            n2661____DOLLAR__6632;
wire            n2662____DOLLAR__6633;
wire            n2663____DOLLAR__6634;
wire            n2664____DOLLAR__6635;
wire            n2665____DOLLAR__6636;
wire            n2666____DOLLAR__6637;
wire            n2667____DOLLAR__6638;
wire            n2668____DOLLAR__6639;
wire            n2669____DOLLAR__6640;
wire            n266____DOLLAR__1029;
wire            n2670____DOLLAR__6641;
wire            n2671____DOLLAR__6642;
wire            n2672____DOLLAR__6643;
wire            n2673____DOLLAR__6644;
wire            n2674____DOLLAR__6645;
wire            n2675____DOLLAR__6646;
wire            n2676____DOLLAR__6647;
wire            n2677____DOLLAR__6648;
wire            n2678____DOLLAR__6649;
wire            n2679____DOLLAR__6650;
wire            n267____DOLLAR__1030;
wire            n2680____DOLLAR__6651;
wire            n2681____DOLLAR__6652;
wire            n2682____DOLLAR__6653;
wire            n2683____DOLLAR__6654;
wire            n2684____DOLLAR__6655;
wire            n2685____DOLLAR__6656;
wire            n2686____DOLLAR__6657;
wire            n2687____DOLLAR__6658;
wire            n2688____DOLLAR__6659;
wire            n2689____DOLLAR__6660;
wire            n268____DOLLAR__1031;
wire            n2690____DOLLAR__6661;
wire            n2691____DOLLAR__6662;
wire            n2692____DOLLAR__6663;
wire            n2693____DOLLAR__6664;
wire            n2694____DOLLAR__6665;
wire            n2695____DOLLAR__6666;
wire            n2696____DOLLAR__6667;
wire            n2697____DOLLAR__6668;
wire            n2698____DOLLAR__6669;
wire            n2699____DOLLAR__6670;
wire            n269____DOLLAR__1032;
wire            n26____DOLLAR__173;
wire            n2700____DOLLAR__6671;
wire            n2701____DOLLAR__6672;
wire            n2702____DOLLAR__6673;
wire            n2703____DOLLAR__6674;
wire            n2704____DOLLAR__6675;
wire            n2705____DOLLAR__6676;
wire            n2706____DOLLAR__6677;
wire            n2707____DOLLAR__6678;
wire            n2708____DOLLAR__6679;
wire            n2709____DOLLAR__6680;
wire            n270____DOLLAR__1033;
wire            n2710____DOLLAR__6681;
wire            n2711____DOLLAR__6682;
wire            n2712____DOLLAR__6683;
wire            n2713____DOLLAR__6684;
wire            n2714____DOLLAR__6685;
wire            n2715____DOLLAR__6686;
wire            n2716____DOLLAR__6687;
wire            n2717____DOLLAR__6688;
wire            n2718____DOLLAR__6689;
wire            n2719____DOLLAR__6690;
wire            n271____DOLLAR__1034;
wire            n2720____DOLLAR__6691;
wire            n2721____DOLLAR__6692;
wire            n2722____DOLLAR__6693;
wire            n2723____DOLLAR__6694;
wire            n2724____DOLLAR__6695;
wire            n2725____DOLLAR__6696;
wire            n2726____DOLLAR__6697;
wire            n2727____DOLLAR__6698;
wire            n2728____DOLLAR__6699;
wire            n2729____DOLLAR__6700;
wire            n272____DOLLAR__1035;
wire            n2730____DOLLAR__6701;
wire            n2731____DOLLAR__6702;
wire            n2732____DOLLAR__6703;
wire            n2733____DOLLAR__6704;
wire            n2734____DOLLAR__6705;
wire            n2735____DOLLAR__6706;
wire            n2736____DOLLAR__6707;
wire            n2737____DOLLAR__6708;
wire            n2738____DOLLAR__6709;
wire            n2739____DOLLAR__6710;
wire            n273____DOLLAR__1036;
wire            n2740____DOLLAR__6711;
wire            n2741____DOLLAR__6712;
wire            n2742____DOLLAR__6713;
wire            n2743____DOLLAR__6714;
wire            n2744____DOLLAR__6715;
wire            n2745____DOLLAR__6716;
wire            n2746____DOLLAR__6717;
wire            n2747____DOLLAR__6718;
wire            n2748____DOLLAR__6719;
wire            n2749____DOLLAR__6720;
wire            n274____DOLLAR__1037;
wire            n2750____DOLLAR__6721;
wire            n2751____DOLLAR__6722;
wire            n2752____DOLLAR__6723;
wire            n2753____DOLLAR__6724;
wire            n2754____DOLLAR__6725;
wire            n2755____DOLLAR__6726;
wire            n2756____DOLLAR__6727;
wire            n2757____DOLLAR__6728;
wire            n2758____DOLLAR__6729;
wire            n2759____DOLLAR__6730;
wire            n275____DOLLAR__1038;
wire            n2760____DOLLAR__6731;
wire            n2761____DOLLAR__6732;
wire            n2762____DOLLAR__6733;
wire            n2763____DOLLAR__6734;
wire            n2764____DOLLAR__6735;
wire            n2765____DOLLAR__6736;
wire            n2766____DOLLAR__6737;
wire            n2767____DOLLAR__6738;
wire            n2768____DOLLAR__6739;
wire            n2769____DOLLAR__6740;
wire            n276____DOLLAR__1039;
wire            n2770____DOLLAR__6741;
wire            n2771____DOLLAR__6742;
wire            n2772____DOLLAR__6743;
wire            n2773____DOLLAR__6744;
wire            n2774____DOLLAR__6745;
wire            n2775____DOLLAR__6746;
wire            n2776____DOLLAR__6747;
wire            n2777____DOLLAR__6748;
wire            n2778____DOLLAR__6749;
wire            n2779____DOLLAR__6750;
wire            n277____DOLLAR__1040;
wire            n2780____DOLLAR__6751;
wire            n2781____DOLLAR__6752;
wire            n2782____DOLLAR__6753;
wire            n2783____DOLLAR__6754;
wire            n2784____DOLLAR__6755;
wire            n2785____DOLLAR__6756;
wire            n2786____DOLLAR__6757;
wire            n2787____DOLLAR__6758;
wire            n2788____DOLLAR__6759;
wire            n2789____DOLLAR__6760;
wire            n278____DOLLAR__1041;
wire            n2790____DOLLAR__6761;
wire            n2791____DOLLAR__6762;
wire            n2792____DOLLAR__6763;
wire            n2793____DOLLAR__6764;
wire            n2794____DOLLAR__6765;
wire            n2795____DOLLAR__6766;
wire            n2796____DOLLAR__6767;
wire     [15:0] n2797____DOLLAR__6770;
wire     [15:0] n2798____DOLLAR__6771;
wire     [15:0] n2799____DOLLAR__6772;
wire            n279____DOLLAR__1042;
wire            n27____DOLLAR__177;
wire     [15:0] n2800____DOLLAR__6773;
wire            n2801____DOLLAR__6778;
wire            n2802____DOLLAR__6782;
wire            n2803____DOLLAR__6786;
wire            n2804____DOLLAR__6788;
wire            n2805____DOLLAR__6789;
wire            n2806____DOLLAR__6794;
wire            n2807____DOLLAR__6798;
wire            n2808____DOLLAR__6802;
wire            n2809____DOLLAR__6806;
wire            n280____DOLLAR__1043;
wire            n2810____DOLLAR__6810;
wire            n2811____DOLLAR__6814;
wire            n2812____DOLLAR__6818;
wire            n2813____DOLLAR__6822;
wire            n2814____DOLLAR__6826;
wire            n2815____DOLLAR__6830;
wire            n2816____DOLLAR__6834;
wire            n2817____DOLLAR__6838;
wire            n2818____DOLLAR__6842;
wire            n2819____DOLLAR__6846;
wire            n281____DOLLAR__1044;
wire            n2820____DOLLAR__6850;
wire            n2821____DOLLAR__6854;
wire            n2822____DOLLAR__6858;
wire            n2823____DOLLAR__6862;
wire            n2824____DOLLAR__6866;
wire            n2825____DOLLAR__6870;
wire            n2826____DOLLAR__6874;
wire            n2827____DOLLAR__6878;
wire            n2828____DOLLAR__6882;
wire            n2829____DOLLAR__6886;
wire            n282____DOLLAR__1045;
wire            n2830____DOLLAR__6890;
wire            n2831____DOLLAR__6894;
wire            n2832____DOLLAR__6898;
wire            n2833____DOLLAR__6902;
wire            n2834____DOLLAR__6906;
wire            n2835____DOLLAR__6910;
wire            n2836____DOLLAR__6914;
wire            n2837____DOLLAR__6918;
wire            n2838____DOLLAR__6922;
wire            n2839____DOLLAR__6926;
wire            n283____DOLLAR__1046;
wire            n2840____DOLLAR__6930;
wire            n2841____DOLLAR__6934;
wire            n2842____DOLLAR__6938;
wire            n2843____DOLLAR__6942;
wire            n2844____DOLLAR__6946;
wire            n2845____DOLLAR__6950;
wire            n2846____DOLLAR__6954;
wire            n2847____DOLLAR__6958;
wire            n2848____DOLLAR__6962;
wire            n2849____DOLLAR__6966;
wire            n284____DOLLAR__1047;
wire            n2850____DOLLAR__6970;
wire            n2851____DOLLAR__6974;
wire            n2852____DOLLAR__6978;
wire            n2853____DOLLAR__6982;
wire            n2854____DOLLAR__6986;
wire            n2855____DOLLAR__6990;
wire            n2856____DOLLAR__6994;
wire            n2857____DOLLAR__6998;
wire            n2858____DOLLAR__7002;
wire            n2859____DOLLAR__7006;
wire            n285____DOLLAR__1048;
wire            n2860____DOLLAR__7010;
wire            n2861____DOLLAR__7014;
wire            n2862____DOLLAR__7018;
wire            n2863____DOLLAR__7022;
wire            n2864____DOLLAR__7026;
wire            n2865____DOLLAR__7030;
wire            n2866____DOLLAR__7034;
wire            n2867____DOLLAR__7038;
wire            n2868____DOLLAR__7042;
wire            n2869____DOLLAR__7046;
wire            n286____DOLLAR__1049;
wire            n2870____DOLLAR__7050;
wire            n2871____DOLLAR__7054;
wire            n2872____DOLLAR__7058;
wire            n2873____DOLLAR__7062;
wire            n2874____DOLLAR__7066;
wire            n2875____DOLLAR__7070;
wire            n2876____DOLLAR__7074;
wire            n2877____DOLLAR__7078;
wire            n2878____DOLLAR__7082;
wire            n2879____DOLLAR__7086;
wire            n287____DOLLAR__1050;
wire            n2880____DOLLAR__7090;
wire            n2881____DOLLAR__7094;
wire            n2882____DOLLAR__7098;
wire            n2883____DOLLAR__7102;
wire            n2884____DOLLAR__7106;
wire            n2885____DOLLAR__7110;
wire            n2886____DOLLAR__7114;
wire            n2887____DOLLAR__7118;
wire            n2888____DOLLAR__7122;
wire            n2889____DOLLAR__7126;
wire            n288____DOLLAR__1051;
wire            n2890____DOLLAR__7130;
wire            n2891____DOLLAR__7134;
wire            n2892____DOLLAR__7138;
wire            n2893____DOLLAR__7142;
wire            n2894____DOLLAR__7146;
wire            n2895____DOLLAR__7150;
wire            n2896____DOLLAR__7154;
wire            n2897____DOLLAR__7158;
wire            n2898____DOLLAR__7162;
wire            n2899____DOLLAR__7166;
wire            n289____DOLLAR__1052;
wire            n28____DOLLAR__181;
wire            n2900____DOLLAR__7170;
wire            n2901____DOLLAR__7174;
wire            n2902____DOLLAR__7178;
wire            n2903____DOLLAR__7182;
wire            n2904____DOLLAR__7186;
wire            n2905____DOLLAR__7190;
wire            n2906____DOLLAR__7194;
wire            n2907____DOLLAR__7198;
wire            n2908____DOLLAR__7202;
wire            n2909____DOLLAR__7206;
wire            n290____DOLLAR__1053;
wire            n2910____DOLLAR__7210;
wire            n2911____DOLLAR__7214;
wire            n2912____DOLLAR__7218;
wire            n2913____DOLLAR__7222;
wire            n2914____DOLLAR__7226;
wire            n2915____DOLLAR__7230;
wire            n2916____DOLLAR__7234;
wire            n2917____DOLLAR__7238;
wire            n2918____DOLLAR__7242;
wire            n2919____DOLLAR__7246;
wire            n291____DOLLAR__1054;
wire            n2920____DOLLAR__7250;
wire            n2921____DOLLAR__7254;
wire            n2922____DOLLAR__7258;
wire            n2923____DOLLAR__7262;
wire            n2924____DOLLAR__7266;
wire            n2925____DOLLAR__7270;
wire            n2926____DOLLAR__7274;
wire            n2927____DOLLAR__7278;
wire            n2928____DOLLAR__7282;
wire            n2929____DOLLAR__7286;
wire            n292____DOLLAR__1055;
wire            n2930____DOLLAR__7290;
wire            n2931____DOLLAR__7294;
wire            n2932____DOLLAR__7298;
wire            n2933____DOLLAR__7302;
wire            n2934____DOLLAR__7306;
wire            n2935____DOLLAR__7310;
wire            n2936____DOLLAR__7314;
wire            n2937____DOLLAR__7318;
wire            n2938____DOLLAR__7322;
wire            n2939____DOLLAR__7326;
wire            n293____DOLLAR__1056;
wire            n2940____DOLLAR__7330;
wire            n2941____DOLLAR__7334;
wire            n2942____DOLLAR__7338;
wire            n2943____DOLLAR__7342;
wire            n2944____DOLLAR__7346;
wire            n2945____DOLLAR__7350;
wire            n2946____DOLLAR__7354;
wire            n2947____DOLLAR__7358;
wire            n2948____DOLLAR__7362;
wire            n2949____DOLLAR__7366;
wire            n294____DOLLAR__1057;
wire            n2950____DOLLAR__7370;
wire            n2951____DOLLAR__7374;
wire            n2952____DOLLAR__7378;
wire            n2953____DOLLAR__7382;
wire            n2954____DOLLAR__7386;
wire            n2955____DOLLAR__7390;
wire            n2956____DOLLAR__7394;
wire            n2957____DOLLAR__7398;
wire            n2958____DOLLAR__7402;
wire            n2959____DOLLAR__7406;
wire            n295____DOLLAR__1058;
wire            n2960____DOLLAR__7410;
wire            n2961____DOLLAR__7414;
wire            n2962____DOLLAR__7418;
wire            n2963____DOLLAR__7422;
wire            n2964____DOLLAR__7426;
wire            n2965____DOLLAR__7430;
wire            n2966____DOLLAR__7434;
wire            n2967____DOLLAR__7438;
wire            n2968____DOLLAR__7442;
wire            n2969____DOLLAR__7446;
wire            n296____DOLLAR__1059;
wire            n2970____DOLLAR__7450;
wire            n2971____DOLLAR__7454;
wire            n2972____DOLLAR__7458;
wire            n2973____DOLLAR__7462;
wire            n2974____DOLLAR__7466;
wire            n2975____DOLLAR__7470;
wire            n2976____DOLLAR__7474;
wire            n2977____DOLLAR__7478;
wire            n2978____DOLLAR__7482;
wire            n2979____DOLLAR__7486;
wire            n297____DOLLAR__1060;
wire            n2980____DOLLAR__7490;
wire            n2981____DOLLAR__7494;
wire            n2982____DOLLAR__7498;
wire            n2983____DOLLAR__7502;
wire            n2984____DOLLAR__7506;
wire            n2985____DOLLAR__7510;
wire            n2986____DOLLAR__7514;
wire            n2987____DOLLAR__7518;
wire            n2988____DOLLAR__7522;
wire            n2989____DOLLAR__7526;
wire            n298____DOLLAR__1061;
wire            n2990____DOLLAR__7530;
wire            n2991____DOLLAR__7534;
wire            n2992____DOLLAR__7538;
wire            n2993____DOLLAR__7542;
wire            n2994____DOLLAR__7546;
wire            n2995____DOLLAR__7550;
wire            n2996____DOLLAR__7554;
wire            n2997____DOLLAR__7558;
wire            n2998____DOLLAR__7562;
wire            n2999____DOLLAR__7566;
wire            n299____DOLLAR__1062;
wire            n29____DOLLAR__185;
wire            n2____DOLLAR__77;
wire            n3000____DOLLAR__7570;
wire            n3001____DOLLAR__7574;
wire            n3002____DOLLAR__7578;
wire            n3003____DOLLAR__7582;
wire            n3004____DOLLAR__7586;
wire            n3005____DOLLAR__7590;
wire            n3006____DOLLAR__7594;
wire            n3007____DOLLAR__7598;
wire            n3008____DOLLAR__7602;
wire            n3009____DOLLAR__7606;
wire            n300____DOLLAR__1063;
wire            n3010____DOLLAR__7610;
wire            n3011____DOLLAR__7614;
wire            n3012____DOLLAR__7618;
wire            n3013____DOLLAR__7622;
wire            n3014____DOLLAR__7626;
wire            n3015____DOLLAR__7630;
wire            n3016____DOLLAR__7634;
wire            n3017____DOLLAR__7638;
wire            n3018____DOLLAR__7642;
wire            n3019____DOLLAR__7646;
wire            n301____DOLLAR__1064;
wire            n3020____DOLLAR__7650;
wire            n3021____DOLLAR__7654;
wire            n3022____DOLLAR__7658;
wire            n3023____DOLLAR__7662;
wire            n3024____DOLLAR__7666;
wire            n3025____DOLLAR__7670;
wire            n3026____DOLLAR__7674;
wire            n3027____DOLLAR__7678;
wire            n3028____DOLLAR__7682;
wire            n3029____DOLLAR__7686;
wire            n302____DOLLAR__1065;
wire            n3030____DOLLAR__7690;
wire            n3031____DOLLAR__7694;
wire            n3032____DOLLAR__7698;
wire            n3033____DOLLAR__7702;
wire            n3034____DOLLAR__7706;
wire            n3035____DOLLAR__7710;
wire            n3036____DOLLAR__7714;
wire            n3037____DOLLAR__7718;
wire            n3038____DOLLAR__7722;
wire            n3039____DOLLAR__7726;
wire            n303____DOLLAR__1066;
wire            n3040____DOLLAR__7730;
wire            n3041____DOLLAR__7734;
wire            n3042____DOLLAR__7738;
wire            n3043____DOLLAR__7742;
wire            n3044____DOLLAR__7746;
wire            n3045____DOLLAR__7750;
wire            n3046____DOLLAR__7754;
wire            n3047____DOLLAR__7758;
wire            n3048____DOLLAR__7762;
wire            n3049____DOLLAR__7766;
wire            n304____DOLLAR__1067;
wire            n3050____DOLLAR__7770;
wire            n3051____DOLLAR__7774;
wire            n3052____DOLLAR__7778;
wire            n3053____DOLLAR__7782;
wire            n3054____DOLLAR__7786;
wire            n3055____DOLLAR__7790;
wire            n3056____DOLLAR__7794;
wire            n3057____DOLLAR__7798;
wire            n3058____DOLLAR__7800;
wire            n3059____DOLLAR__7802;
wire            n305____DOLLAR__1068;
wire            n3060____DOLLAR__7803;
wire            n3061____DOLLAR__7804;
wire            n3062____DOLLAR__7805;
wire            n3063____DOLLAR__7806;
wire            n3064____DOLLAR__7807;
wire            n3065____DOLLAR__7808;
wire            n3066____DOLLAR__7809;
wire            n3067____DOLLAR__7810;
wire            n3068____DOLLAR__7811;
wire            n3069____DOLLAR__7812;
wire            n306____DOLLAR__1069;
wire            n3070____DOLLAR__7813;
wire            n3071____DOLLAR__7814;
wire            n3072____DOLLAR__7815;
wire            n3073____DOLLAR__7816;
wire            n3074____DOLLAR__7817;
wire            n3075____DOLLAR__7818;
wire            n3076____DOLLAR__7819;
wire            n3077____DOLLAR__7820;
wire            n3078____DOLLAR__7821;
wire            n3079____DOLLAR__7822;
wire            n307____DOLLAR__1070;
wire            n3080____DOLLAR__7823;
wire            n3081____DOLLAR__7824;
wire            n3082____DOLLAR__7825;
wire            n3083____DOLLAR__7826;
wire            n3084____DOLLAR__7827;
wire            n3085____DOLLAR__7828;
wire            n3086____DOLLAR__7829;
wire            n3087____DOLLAR__7830;
wire            n3088____DOLLAR__7831;
wire            n3089____DOLLAR__7832;
wire            n308____DOLLAR__1071;
wire            n3090____DOLLAR__7833;
wire            n3091____DOLLAR__7834;
wire            n3092____DOLLAR__7835;
wire            n3093____DOLLAR__7836;
wire            n3094____DOLLAR__7837;
wire            n3095____DOLLAR__7838;
wire            n3096____DOLLAR__7839;
wire            n3097____DOLLAR__7840;
wire            n3098____DOLLAR__7841;
wire            n3099____DOLLAR__7842;
wire            n309____DOLLAR__1072;
wire            n30____DOLLAR__189;
wire            n3100____DOLLAR__7843;
wire            n3101____DOLLAR__7844;
wire            n3102____DOLLAR__7845;
wire            n3103____DOLLAR__7846;
wire            n3104____DOLLAR__7847;
wire            n3105____DOLLAR__7848;
wire            n3106____DOLLAR__7849;
wire            n3107____DOLLAR__7850;
wire            n3108____DOLLAR__7851;
wire            n3109____DOLLAR__7852;
wire            n310____DOLLAR__1073;
wire            n3110____DOLLAR__7853;
wire            n3111____DOLLAR__7854;
wire            n3112____DOLLAR__7855;
wire            n3113____DOLLAR__7856;
wire            n3114____DOLLAR__7857;
wire            n3115____DOLLAR__7858;
wire            n3116____DOLLAR__7859;
wire            n3117____DOLLAR__7860;
wire            n3118____DOLLAR__7861;
wire            n3119____DOLLAR__7862;
wire            n311____DOLLAR__1074;
wire            n3120____DOLLAR__7863;
wire            n3121____DOLLAR__7864;
wire            n3122____DOLLAR__7865;
wire            n3123____DOLLAR__7866;
wire            n3124____DOLLAR__7867;
wire            n3125____DOLLAR__7868;
wire            n3126____DOLLAR__7869;
wire            n3127____DOLLAR__7870;
wire            n3128____DOLLAR__7871;
wire            n3129____DOLLAR__7872;
wire            n312____DOLLAR__1075;
wire            n3130____DOLLAR__7873;
wire            n3131____DOLLAR__7874;
wire            n3132____DOLLAR__7875;
wire            n3133____DOLLAR__7876;
wire            n3134____DOLLAR__7877;
wire            n3135____DOLLAR__7878;
wire            n3136____DOLLAR__7879;
wire            n3137____DOLLAR__7880;
wire            n3138____DOLLAR__7881;
wire            n3139____DOLLAR__7882;
wire            n313____DOLLAR__1076;
wire            n3140____DOLLAR__7883;
wire            n3141____DOLLAR__7884;
wire            n3142____DOLLAR__7885;
wire            n3143____DOLLAR__7886;
wire            n3144____DOLLAR__7887;
wire            n3145____DOLLAR__7888;
wire            n3146____DOLLAR__7889;
wire            n3147____DOLLAR__7890;
wire            n3148____DOLLAR__7891;
wire            n3149____DOLLAR__7892;
wire            n314____DOLLAR__1077;
wire            n3150____DOLLAR__7893;
wire            n3151____DOLLAR__7894;
wire            n3152____DOLLAR__7895;
wire            n3153____DOLLAR__7896;
wire            n3154____DOLLAR__7897;
wire            n3155____DOLLAR__7898;
wire            n3156____DOLLAR__7899;
wire            n3157____DOLLAR__7900;
wire            n3158____DOLLAR__7901;
wire            n3159____DOLLAR__7902;
wire            n315____DOLLAR__1078;
wire            n3160____DOLLAR__7903;
wire            n3161____DOLLAR__7904;
wire            n3162____DOLLAR__7905;
wire            n3163____DOLLAR__7906;
wire            n3164____DOLLAR__7907;
wire            n3165____DOLLAR__7908;
wire            n3166____DOLLAR__7909;
wire            n3167____DOLLAR__7910;
wire            n3168____DOLLAR__7911;
wire            n3169____DOLLAR__7912;
wire            n316____DOLLAR__1079;
wire            n3170____DOLLAR__7913;
wire            n3171____DOLLAR__7914;
wire            n3172____DOLLAR__7915;
wire            n3173____DOLLAR__7916;
wire            n3174____DOLLAR__7917;
wire            n3175____DOLLAR__7918;
wire            n3176____DOLLAR__7919;
wire            n3177____DOLLAR__7920;
wire            n3178____DOLLAR__7921;
wire            n3179____DOLLAR__7922;
wire            n317____DOLLAR__1080;
wire            n3180____DOLLAR__7923;
wire            n3181____DOLLAR__7924;
wire            n3182____DOLLAR__7925;
wire            n3183____DOLLAR__7926;
wire            n3184____DOLLAR__7927;
wire            n3185____DOLLAR__7928;
wire            n3186____DOLLAR__7929;
wire            n3187____DOLLAR__7930;
wire            n3188____DOLLAR__7931;
wire            n3189____DOLLAR__7932;
wire            n318____DOLLAR__1081;
wire            n3190____DOLLAR__7933;
wire            n3191____DOLLAR__7934;
wire            n3192____DOLLAR__7935;
wire            n3193____DOLLAR__7936;
wire            n3194____DOLLAR__7937;
wire            n3195____DOLLAR__7938;
wire            n3196____DOLLAR__7939;
wire            n3197____DOLLAR__7940;
wire            n3198____DOLLAR__7941;
wire            n3199____DOLLAR__7942;
wire            n319____DOLLAR__1082;
wire            n31____DOLLAR__193;
wire            n3200____DOLLAR__7943;
wire            n3201____DOLLAR__7944;
wire            n3202____DOLLAR__7945;
wire            n3203____DOLLAR__7946;
wire            n3204____DOLLAR__7947;
wire            n3205____DOLLAR__7948;
wire            n3206____DOLLAR__7949;
wire            n3207____DOLLAR__7950;
wire            n3208____DOLLAR__7951;
wire            n3209____DOLLAR__7952;
wire            n320____DOLLAR__1083;
wire            n3210____DOLLAR__7953;
wire            n3211____DOLLAR__7954;
wire            n3212____DOLLAR__7955;
wire            n3213____DOLLAR__7956;
wire            n3214____DOLLAR__7957;
wire            n3215____DOLLAR__7958;
wire            n3216____DOLLAR__7959;
wire            n3217____DOLLAR__7960;
wire            n3218____DOLLAR__7961;
wire            n3219____DOLLAR__7962;
wire            n321____DOLLAR__1084;
wire            n3220____DOLLAR__7963;
wire            n3221____DOLLAR__7964;
wire            n3222____DOLLAR__7965;
wire            n3223____DOLLAR__7966;
wire            n3224____DOLLAR__7967;
wire            n3225____DOLLAR__7968;
wire            n3226____DOLLAR__7969;
wire            n3227____DOLLAR__7970;
wire            n3228____DOLLAR__7971;
wire            n3229____DOLLAR__7972;
wire            n322____DOLLAR__1085;
wire            n3230____DOLLAR__7973;
wire            n3231____DOLLAR__7974;
wire            n3232____DOLLAR__7975;
wire            n3233____DOLLAR__7976;
wire            n3234____DOLLAR__7977;
wire            n3235____DOLLAR__7978;
wire            n3236____DOLLAR__7979;
wire            n3237____DOLLAR__7980;
wire            n3238____DOLLAR__7981;
wire            n3239____DOLLAR__7982;
wire            n323____DOLLAR__1086;
wire            n3240____DOLLAR__7983;
wire            n3241____DOLLAR__7984;
wire            n3242____DOLLAR__7985;
wire            n3243____DOLLAR__7986;
wire            n3244____DOLLAR__7987;
wire            n3245____DOLLAR__7988;
wire            n3246____DOLLAR__7989;
wire            n3247____DOLLAR__7990;
wire            n3248____DOLLAR__7991;
wire            n3249____DOLLAR__7992;
wire            n324____DOLLAR__1087;
wire            n3250____DOLLAR__7993;
wire            n3251____DOLLAR__7994;
wire            n3252____DOLLAR__7995;
wire            n3253____DOLLAR__7996;
wire            n3254____DOLLAR__7997;
wire            n3255____DOLLAR__7998;
wire            n3256____DOLLAR__7999;
wire            n3257____DOLLAR__8000;
wire            n3258____DOLLAR__8001;
wire            n3259____DOLLAR__8002;
wire            n325____DOLLAR__1088;
wire            n3260____DOLLAR__8003;
wire            n3261____DOLLAR__8004;
wire            n3262____DOLLAR__8005;
wire            n3263____DOLLAR__8006;
wire            n3264____DOLLAR__8007;
wire            n3265____DOLLAR__8008;
wire            n3266____DOLLAR__8009;
wire            n3267____DOLLAR__8010;
wire            n3268____DOLLAR__8011;
wire            n3269____DOLLAR__8012;
wire            n326____DOLLAR__1089;
wire            n3270____DOLLAR__8013;
wire            n3271____DOLLAR__8014;
wire            n3272____DOLLAR__8015;
wire            n3273____DOLLAR__8016;
wire            n3274____DOLLAR__8017;
wire            n3275____DOLLAR__8018;
wire            n3276____DOLLAR__8019;
wire            n3277____DOLLAR__8020;
wire            n3278____DOLLAR__8021;
wire            n3279____DOLLAR__8022;
wire            n327____DOLLAR__1090;
wire            n3280____DOLLAR__8023;
wire            n3281____DOLLAR__8024;
wire            n3282____DOLLAR__8025;
wire            n3283____DOLLAR__8026;
wire            n3284____DOLLAR__8027;
wire            n3285____DOLLAR__8028;
wire            n3286____DOLLAR__8029;
wire            n3287____DOLLAR__8030;
wire            n3288____DOLLAR__8031;
wire            n3289____DOLLAR__8032;
wire            n328____DOLLAR__1091;
wire            n3290____DOLLAR__8033;
wire            n3291____DOLLAR__8034;
wire            n3292____DOLLAR__8035;
wire            n3293____DOLLAR__8036;
wire            n3294____DOLLAR__8037;
wire            n3295____DOLLAR__8038;
wire            n3296____DOLLAR__8039;
wire            n3297____DOLLAR__8040;
wire            n3298____DOLLAR__8041;
wire            n3299____DOLLAR__8042;
wire            n329____DOLLAR__1092;
wire            n32____DOLLAR__197;
wire            n3300____DOLLAR__8043;
wire            n3301____DOLLAR__8044;
wire            n3302____DOLLAR__8045;
wire            n3303____DOLLAR__8046;
wire            n3304____DOLLAR__8047;
wire            n3305____DOLLAR__8048;
wire            n3306____DOLLAR__8049;
wire            n3307____DOLLAR__8050;
wire            n3308____DOLLAR__8051;
wire            n3309____DOLLAR__8052;
wire            n330____DOLLAR__1093;
wire            n3310____DOLLAR__8053;
wire      [7:0] n3311____DOLLAR__8056;
wire      [7:0] n3312____DOLLAR__8057;
wire     [15:0] n3313____DOLLAR__203215;
wire     [15:0] n3314____DOLLAR__203218;
wire            n3315____DOLLAR__203842;
wire            n3316____DOLLAR__204105;
wire            n3317____DOLLAR__204106;
wire            n3318____DOLLAR__204104;
wire     [15:0] n3319____DOLLAR__203240;
wire            n331____DOLLAR__1094;
wire            n3320____DOLLAR__203836;
wire            n3321____DOLLAR__203829;
wire            n3322____DOLLAR__203831;
wire            n3323____DOLLAR__203833;
wire            n3324____DOLLAR__203838;
wire            n3325____DOLLAR__204108;
wire            n3326____DOLLAR__204109;
wire            n3327____DOLLAR__204107;
wire            n3328____DOLLAR__203301;
wire            n3329____DOLLAR__203296;
wire            n332____DOLLAR__1095;
wire      [7:0] n3330____DOLLAR__203286;
wire     [15:0] n3331____DOLLAR__203292;
wire            n3332____DOLLAR__203283;
wire      [7:0] n3333____DOLLAR__203273;
wire     [15:0] n3334____DOLLAR__203279;
wire     [15:0] n3335____DOLLAR__203285;
wire     [15:0] n3336____DOLLAR__203298;
wire     [15:0] n3337____DOLLAR__203303;
wire            n3338____DOLLAR__203270;
wire            n3339____DOLLAR__203265;
wire            n333____DOLLAR__1096;
wire      [7:0] n3340____DOLLAR__203255;
wire     [15:0] n3341____DOLLAR__203261;
wire            n3342____DOLLAR__203252;
wire      [7:0] n3343____DOLLAR__203242;
wire     [15:0] n3344____DOLLAR__203248;
wire     [15:0] n3345____DOLLAR__203254;
wire     [15:0] n3346____DOLLAR__203267;
wire     [15:0] n3347____DOLLAR__203272;
wire            n3348____DOLLAR__203556;
wire     [15:0] n3349____DOLLAR__203542;
wire            n334____DOLLAR__1097;
wire            n3350____DOLLAR__203545;
wire      [7:0] n3351____DOLLAR__203538;
wire      [7:0] n3352____DOLLAR__203547;
wire     [15:0] n3353____DOLLAR__203526;
wire            n3354____DOLLAR__203529;
wire      [7:0] n3355____DOLLAR__203522;
wire      [7:0] n3356____DOLLAR__203531;
wire     [15:0] n3357____DOLLAR__203510;
wire            n3358____DOLLAR__203513;
wire      [7:0] n3359____DOLLAR__203506;
wire            n335____DOLLAR__1098;
wire      [7:0] n3360____DOLLAR__203515;
wire     [15:0] n3361____DOLLAR__203494;
wire            n3362____DOLLAR__203497;
wire      [7:0] n3363____DOLLAR__203490;
wire      [7:0] n3364____DOLLAR__203499;
wire     [15:0] n3365____DOLLAR__203478;
wire            n3366____DOLLAR__203481;
wire      [7:0] n3367____DOLLAR__203474;
wire      [7:0] n3368____DOLLAR__203483;
wire     [15:0] n3369____DOLLAR__203462;
wire            n336____DOLLAR__1099;
wire            n3370____DOLLAR__203465;
wire      [7:0] n3371____DOLLAR__203458;
wire      [7:0] n3372____DOLLAR__203467;
wire     [15:0] n3373____DOLLAR__203446;
wire            n3374____DOLLAR__203449;
wire      [7:0] n3375____DOLLAR__203442;
wire      [7:0] n3376____DOLLAR__203451;
wire     [15:0] n3377____DOLLAR__203430;
wire            n3378____DOLLAR__203433;
wire      [7:0] n3379____DOLLAR__203426;
wire            n337____DOLLAR__1100;
wire      [7:0] n3380____DOLLAR__203435;
wire     [15:0] n3381____DOLLAR__203414;
wire            n3382____DOLLAR__203417;
wire      [7:0] n3383____DOLLAR__203410;
wire      [7:0] n3384____DOLLAR__203419;
wire     [15:0] n3385____DOLLAR__203398;
wire            n3386____DOLLAR__203401;
wire      [7:0] n3387____DOLLAR__203394;
wire      [7:0] n3388____DOLLAR__203403;
wire     [15:0] n3389____DOLLAR__203382;
wire            n338____DOLLAR__1101;
wire            n3390____DOLLAR__203385;
wire      [7:0] n3391____DOLLAR__203378;
wire      [7:0] n3392____DOLLAR__203387;
wire     [15:0] n3393____DOLLAR__203366;
wire            n3394____DOLLAR__203369;
wire      [7:0] n3395____DOLLAR__203362;
wire      [7:0] n3396____DOLLAR__203371;
wire     [15:0] n3397____DOLLAR__203350;
wire            n3398____DOLLAR__203353;
wire      [7:0] n3399____DOLLAR__203346;
wire            n339____DOLLAR__1102;
wire            n33____DOLLAR__201;
wire      [7:0] n3400____DOLLAR__203355;
wire     [15:0] n3401____DOLLAR__203334;
wire            n3402____DOLLAR__203337;
wire      [7:0] n3403____DOLLAR__203330;
wire      [7:0] n3404____DOLLAR__203339;
wire     [15:0] n3405____DOLLAR__203318;
wire            n3406____DOLLAR__203321;
wire      [7:0] n3407____DOLLAR__203314;
wire      [7:0] n3408____DOLLAR__203323;
wire     [15:0] n3409____DOLLAR__203308;
wire            n340____DOLLAR__1103;
wire            n3410____DOLLAR__203311;
wire      [7:0] n3411____DOLLAR__203304;
wire      [7:0] n3412____DOLLAR__203313;
wire     [15:0] n3413____DOLLAR__203328;
wire     [23:0] n3414____DOLLAR__203344;
wire     [31:0] n3415____DOLLAR__203360;
wire     [39:0] n3416____DOLLAR__203376;
wire     [47:0] n3417____DOLLAR__203392;
wire     [55:0] n3418____DOLLAR__203408;
wire     [63:0] n3419____DOLLAR__203424;
wire            n341____DOLLAR__1104;
wire     [71:0] n3420____DOLLAR__203440;
wire     [79:0] n3421____DOLLAR__203456;
wire     [87:0] n3422____DOLLAR__203472;
wire     [95:0] n3423____DOLLAR__203488;
wire    [103:0] n3424____DOLLAR__203504;
wire    [111:0] n3425____DOLLAR__203520;
wire    [119:0] n3426____DOLLAR__203536;
wire    [127:0] n3427____DOLLAR__203552;
wire    [127:0] n3428____DOLLAR__203558;
wire            n3429____DOLLAR__203811;
wire            n342____DOLLAR__1105;
wire     [15:0] n3430____DOLLAR__203797;
wire            n3431____DOLLAR__203800;
wire      [7:0] n3432____DOLLAR__203793;
wire      [7:0] n3433____DOLLAR__203802;
wire     [15:0] n3434____DOLLAR__203781;
wire            n3435____DOLLAR__203784;
wire      [7:0] n3436____DOLLAR__203777;
wire      [7:0] n3437____DOLLAR__203786;
wire     [15:0] n3438____DOLLAR__203765;
wire            n3439____DOLLAR__203768;
wire            n343____DOLLAR__1106;
wire      [7:0] n3440____DOLLAR__203761;
wire      [7:0] n3441____DOLLAR__203770;
wire     [15:0] n3442____DOLLAR__203749;
wire            n3443____DOLLAR__203752;
wire      [7:0] n3444____DOLLAR__203745;
wire      [7:0] n3445____DOLLAR__203754;
wire     [15:0] n3446____DOLLAR__203733;
wire            n3447____DOLLAR__203736;
wire      [7:0] n3448____DOLLAR__203729;
wire      [7:0] n3449____DOLLAR__203738;
wire            n344____DOLLAR__1107;
wire     [15:0] n3450____DOLLAR__203717;
wire            n3451____DOLLAR__203720;
wire      [7:0] n3452____DOLLAR__203713;
wire      [7:0] n3453____DOLLAR__203722;
wire     [15:0] n3454____DOLLAR__203701;
wire            n3455____DOLLAR__203704;
wire      [7:0] n3456____DOLLAR__203697;
wire      [7:0] n3457____DOLLAR__203706;
wire     [15:0] n3458____DOLLAR__203685;
wire            n3459____DOLLAR__203688;
wire            n345____DOLLAR__1108;
wire      [7:0] n3460____DOLLAR__203681;
wire      [7:0] n3461____DOLLAR__203690;
wire     [15:0] n3462____DOLLAR__203669;
wire            n3463____DOLLAR__203672;
wire      [7:0] n3464____DOLLAR__203665;
wire      [7:0] n3465____DOLLAR__203674;
wire     [15:0] n3466____DOLLAR__203653;
wire            n3467____DOLLAR__203656;
wire      [7:0] n3468____DOLLAR__203649;
wire      [7:0] n3469____DOLLAR__203658;
wire            n346____DOLLAR__1109;
wire     [15:0] n3470____DOLLAR__203637;
wire            n3471____DOLLAR__203640;
wire      [7:0] n3472____DOLLAR__203633;
wire      [7:0] n3473____DOLLAR__203642;
wire     [15:0] n3474____DOLLAR__203621;
wire            n3475____DOLLAR__203624;
wire      [7:0] n3476____DOLLAR__203617;
wire      [7:0] n3477____DOLLAR__203626;
wire     [15:0] n3478____DOLLAR__203605;
wire            n3479____DOLLAR__203608;
wire            n347____DOLLAR__1110;
wire      [7:0] n3480____DOLLAR__203601;
wire      [7:0] n3481____DOLLAR__203610;
wire     [15:0] n3482____DOLLAR__203589;
wire            n3483____DOLLAR__203592;
wire      [7:0] n3484____DOLLAR__203585;
wire      [7:0] n3485____DOLLAR__203594;
wire     [15:0] n3486____DOLLAR__203573;
wire            n3487____DOLLAR__203576;
wire      [7:0] n3488____DOLLAR__203569;
wire      [7:0] n3489____DOLLAR__203578;
wire            n348____DOLLAR__1111;
wire     [15:0] n3490____DOLLAR__203563;
wire            n3491____DOLLAR__203566;
wire      [7:0] n3492____DOLLAR__203559;
wire      [7:0] n3493____DOLLAR__203568;
wire     [15:0] n3494____DOLLAR__203583;
wire     [23:0] n3495____DOLLAR__203599;
wire     [31:0] n3496____DOLLAR__203615;
wire     [39:0] n3497____DOLLAR__203631;
wire     [47:0] n3498____DOLLAR__203647;
wire     [55:0] n3499____DOLLAR__203663;
wire            n349____DOLLAR__1112;
wire            n34____DOLLAR__205;
wire     [63:0] n3500____DOLLAR__203679;
wire     [71:0] n3501____DOLLAR__203695;
wire     [79:0] n3502____DOLLAR__203711;
wire     [87:0] n3503____DOLLAR__203727;
wire     [95:0] n3504____DOLLAR__203743;
wire    [103:0] n3505____DOLLAR__203759;
wire    [111:0] n3506____DOLLAR__203775;
wire    [119:0] n3507____DOLLAR__203791;
wire    [127:0] n3508____DOLLAR__203807;
wire    [127:0] n3509____DOLLAR__203813;
wire            n350____DOLLAR__1113;
wire            n3510____DOLLAR__203823;
wire            n3511____DOLLAR__203818;
wire      [1:0] n3512____DOLLAR__203820;
wire      [1:0] n3513____DOLLAR__203825;
wire            n351____DOLLAR__1114;
wire            n352____DOLLAR__1115;
wire            n353____DOLLAR__1116;
wire            n354____DOLLAR__1117;
wire            n355____DOLLAR__1118;
wire            n356____DOLLAR__1119;
wire            n357____DOLLAR__1120;
wire            n358____DOLLAR__1121;
wire            n359____DOLLAR__1122;
wire            n35____DOLLAR__209;
wire            n360____DOLLAR__1123;
wire            n361____DOLLAR__1124;
wire            n362____DOLLAR__1125;
wire            n363____DOLLAR__1126;
wire            n364____DOLLAR__1127;
wire            n365____DOLLAR__1128;
wire            n366____DOLLAR__1129;
wire            n367____DOLLAR__1130;
wire            n368____DOLLAR__1131;
wire            n369____DOLLAR__1132;
wire            n36____DOLLAR__213;
wire            n370____DOLLAR__1133;
wire            n371____DOLLAR__1134;
wire            n372____DOLLAR__1135;
wire            n373____DOLLAR__1136;
wire            n374____DOLLAR__1137;
wire            n375____DOLLAR__1138;
wire            n376____DOLLAR__1139;
wire            n377____DOLLAR__1140;
wire            n378____DOLLAR__1141;
wire            n379____DOLLAR__1142;
wire            n37____DOLLAR__217;
wire            n380____DOLLAR__1143;
wire            n381____DOLLAR__1144;
wire            n382____DOLLAR__1145;
wire            n383____DOLLAR__1146;
wire            n384____DOLLAR__1147;
wire            n385____DOLLAR__1148;
wire            n386____DOLLAR__1149;
wire            n387____DOLLAR__1150;
wire            n388____DOLLAR__1151;
wire            n389____DOLLAR__1152;
wire            n38____DOLLAR__221;
wire            n390____DOLLAR__1153;
wire            n391____DOLLAR__1154;
wire            n392____DOLLAR__1155;
wire            n393____DOLLAR__1156;
wire            n394____DOLLAR__1157;
wire            n395____DOLLAR__1158;
wire            n396____DOLLAR__1159;
wire            n397____DOLLAR__1160;
wire            n398____DOLLAR__1161;
wire            n399____DOLLAR__1162;
wire            n39____DOLLAR__225;
wire            n3____DOLLAR__81;
wire            n400____DOLLAR__1163;
wire            n401____DOLLAR__1164;
wire            n402____DOLLAR__1165;
wire            n403____DOLLAR__1166;
wire            n404____DOLLAR__1167;
wire            n405____DOLLAR__1168;
wire            n406____DOLLAR__1169;
wire            n407____DOLLAR__1170;
wire            n408____DOLLAR__1171;
wire            n409____DOLLAR__1172;
wire            n40____DOLLAR__229;
wire            n410____DOLLAR__1173;
wire            n411____DOLLAR__1174;
wire            n412____DOLLAR__1175;
wire            n413____DOLLAR__1176;
wire            n414____DOLLAR__1177;
wire            n415____DOLLAR__1178;
wire            n416____DOLLAR__1179;
wire            n417____DOLLAR__1180;
wire            n418____DOLLAR__1181;
wire            n419____DOLLAR__1182;
wire            n41____DOLLAR__233;
wire            n420____DOLLAR__1183;
wire            n421____DOLLAR__1184;
wire            n422____DOLLAR__1185;
wire            n423____DOLLAR__1186;
wire            n424____DOLLAR__1187;
wire            n425____DOLLAR__1188;
wire            n426____DOLLAR__1189;
wire            n427____DOLLAR__1190;
wire            n428____DOLLAR__1191;
wire            n429____DOLLAR__1192;
wire            n42____DOLLAR__237;
wire            n430____DOLLAR__1193;
wire            n431____DOLLAR__1194;
wire            n432____DOLLAR__1195;
wire            n433____DOLLAR__1196;
wire            n434____DOLLAR__1197;
wire            n435____DOLLAR__1198;
wire            n436____DOLLAR__1199;
wire            n437____DOLLAR__1200;
wire            n438____DOLLAR__1201;
wire            n439____DOLLAR__1202;
wire            n43____DOLLAR__241;
wire            n440____DOLLAR__1203;
wire            n441____DOLLAR__1204;
wire            n442____DOLLAR__1205;
wire            n443____DOLLAR__1206;
wire            n444____DOLLAR__1207;
wire            n445____DOLLAR__1208;
wire            n446____DOLLAR__1209;
wire            n447____DOLLAR__1210;
wire            n448____DOLLAR__1211;
wire            n449____DOLLAR__1212;
wire            n44____DOLLAR__245;
wire            n450____DOLLAR__1213;
wire            n451____DOLLAR__1214;
wire            n452____DOLLAR__1215;
wire            n453____DOLLAR__1216;
wire            n454____DOLLAR__1217;
wire            n455____DOLLAR__1218;
wire            n456____DOLLAR__1219;
wire            n457____DOLLAR__1220;
wire            n458____DOLLAR__1221;
wire            n459____DOLLAR__1222;
wire            n45____DOLLAR__249;
wire            n460____DOLLAR__1223;
wire     [15:0] n461____DOLLAR__1228;
wire      [7:0] n462____DOLLAR__1230;
wire      [7:0] n463____DOLLAR__1232;
wire            n464____DOLLAR__1237;
wire            n465____DOLLAR__1241;
wire            n466____DOLLAR__1245;
wire            n467____DOLLAR__1249;
wire            n468____DOLLAR__1253;
wire            n469____DOLLAR__1257;
wire            n46____DOLLAR__253;
wire            n470____DOLLAR__1261;
wire            n471____DOLLAR__1265;
wire            n472____DOLLAR__1269;
wire            n473____DOLLAR__1273;
wire            n474____DOLLAR__1277;
wire            n475____DOLLAR__1281;
wire            n476____DOLLAR__1285;
wire            n477____DOLLAR__1289;
wire            n478____DOLLAR__1293;
wire            n479____DOLLAR__1297;
wire            n47____DOLLAR__257;
wire            n480____DOLLAR__1301;
wire            n481____DOLLAR__1305;
wire            n482____DOLLAR__1309;
wire            n483____DOLLAR__1313;
wire            n484____DOLLAR__1317;
wire            n485____DOLLAR__1321;
wire            n486____DOLLAR__1325;
wire            n487____DOLLAR__1329;
wire            n488____DOLLAR__1333;
wire            n489____DOLLAR__1337;
wire            n48____DOLLAR__261;
wire            n490____DOLLAR__1341;
wire            n491____DOLLAR__1345;
wire            n492____DOLLAR__1349;
wire            n493____DOLLAR__1353;
wire            n494____DOLLAR__1357;
wire            n495____DOLLAR__1361;
wire            n496____DOLLAR__1365;
wire            n497____DOLLAR__1369;
wire            n498____DOLLAR__1373;
wire            n499____DOLLAR__1377;
wire            n49____DOLLAR__265;
wire            n4____DOLLAR__85;
wire            n500____DOLLAR__1381;
wire            n501____DOLLAR__1385;
wire            n502____DOLLAR__1389;
wire            n503____DOLLAR__1393;
wire            n504____DOLLAR__1397;
wire            n505____DOLLAR__1401;
wire            n506____DOLLAR__1405;
wire            n507____DOLLAR__1409;
wire            n508____DOLLAR__1413;
wire            n509____DOLLAR__1417;
wire            n50____DOLLAR__269;
wire            n510____DOLLAR__1421;
wire            n511____DOLLAR__1425;
wire            n512____DOLLAR__1429;
wire            n513____DOLLAR__1433;
wire            n514____DOLLAR__1437;
wire            n515____DOLLAR__1441;
wire            n516____DOLLAR__1445;
wire            n517____DOLLAR__1449;
wire            n518____DOLLAR__1453;
wire            n519____DOLLAR__1457;
wire            n51____DOLLAR__273;
wire            n520____DOLLAR__1461;
wire            n521____DOLLAR__1465;
wire            n522____DOLLAR__1469;
wire            n523____DOLLAR__1473;
wire            n524____DOLLAR__1477;
wire            n525____DOLLAR__1481;
wire            n526____DOLLAR__1485;
wire            n527____DOLLAR__1489;
wire            n528____DOLLAR__1493;
wire            n529____DOLLAR__1497;
wire            n52____DOLLAR__277;
wire            n530____DOLLAR__1501;
wire            n531____DOLLAR__1505;
wire            n532____DOLLAR__1509;
wire            n533____DOLLAR__1513;
wire            n534____DOLLAR__1517;
wire            n535____DOLLAR__1521;
wire            n536____DOLLAR__1525;
wire            n537____DOLLAR__1529;
wire            n538____DOLLAR__1533;
wire            n539____DOLLAR__1537;
wire            n53____DOLLAR__281;
wire            n540____DOLLAR__1541;
wire            n541____DOLLAR__1545;
wire            n542____DOLLAR__1549;
wire            n543____DOLLAR__1553;
wire            n544____DOLLAR__1557;
wire            n545____DOLLAR__1561;
wire            n546____DOLLAR__1565;
wire            n547____DOLLAR__1569;
wire            n548____DOLLAR__1573;
wire            n549____DOLLAR__1577;
wire            n54____DOLLAR__285;
wire            n550____DOLLAR__1581;
wire            n551____DOLLAR__1585;
wire            n552____DOLLAR__1589;
wire            n553____DOLLAR__1593;
wire            n554____DOLLAR__1597;
wire            n555____DOLLAR__1601;
wire            n556____DOLLAR__1605;
wire            n557____DOLLAR__1609;
wire            n558____DOLLAR__1613;
wire            n559____DOLLAR__1617;
wire            n55____DOLLAR__289;
wire            n560____DOLLAR__1621;
wire            n561____DOLLAR__1625;
wire            n562____DOLLAR__1629;
wire            n563____DOLLAR__1633;
wire            n564____DOLLAR__1637;
wire            n565____DOLLAR__1641;
wire            n566____DOLLAR__1645;
wire            n567____DOLLAR__1649;
wire            n568____DOLLAR__1653;
wire            n569____DOLLAR__1657;
wire            n56____DOLLAR__293;
wire            n570____DOLLAR__1661;
wire            n571____DOLLAR__1665;
wire            n572____DOLLAR__1669;
wire            n573____DOLLAR__1673;
wire            n574____DOLLAR__1677;
wire            n575____DOLLAR__1681;
wire            n576____DOLLAR__1685;
wire            n577____DOLLAR__1689;
wire            n578____DOLLAR__1693;
wire            n579____DOLLAR__1697;
wire            n57____DOLLAR__297;
wire            n580____DOLLAR__1701;
wire            n581____DOLLAR__1705;
wire            n582____DOLLAR__1709;
wire            n583____DOLLAR__1713;
wire            n584____DOLLAR__1717;
wire            n585____DOLLAR__1721;
wire            n586____DOLLAR__1725;
wire            n587____DOLLAR__1729;
wire            n588____DOLLAR__1733;
wire            n589____DOLLAR__1737;
wire            n58____DOLLAR__301;
wire            n590____DOLLAR__1741;
wire            n591____DOLLAR__1745;
wire            n592____DOLLAR__1749;
wire            n593____DOLLAR__1753;
wire            n594____DOLLAR__1757;
wire            n595____DOLLAR__1761;
wire            n596____DOLLAR__1765;
wire            n597____DOLLAR__1769;
wire            n598____DOLLAR__1773;
wire            n599____DOLLAR__1777;
wire            n59____DOLLAR__305;
wire            n5____DOLLAR__89;
wire            n600____DOLLAR__1781;
wire            n601____DOLLAR__1785;
wire            n602____DOLLAR__1789;
wire            n603____DOLLAR__1793;
wire            n604____DOLLAR__1797;
wire            n605____DOLLAR__1801;
wire            n606____DOLLAR__1805;
wire            n607____DOLLAR__1809;
wire            n608____DOLLAR__1813;
wire            n609____DOLLAR__1817;
wire            n60____DOLLAR__309;
wire            n610____DOLLAR__1821;
wire            n611____DOLLAR__1825;
wire            n612____DOLLAR__1829;
wire            n613____DOLLAR__1833;
wire            n614____DOLLAR__1837;
wire            n615____DOLLAR__1841;
wire            n616____DOLLAR__1845;
wire            n617____DOLLAR__1849;
wire            n618____DOLLAR__1853;
wire            n619____DOLLAR__1857;
wire            n61____DOLLAR__313;
wire            n620____DOLLAR__1861;
wire            n621____DOLLAR__1865;
wire            n622____DOLLAR__1869;
wire            n623____DOLLAR__1873;
wire            n624____DOLLAR__1877;
wire            n625____DOLLAR__1881;
wire            n626____DOLLAR__1885;
wire            n627____DOLLAR__1889;
wire            n628____DOLLAR__1893;
wire            n629____DOLLAR__1897;
wire            n62____DOLLAR__317;
wire            n630____DOLLAR__1901;
wire            n631____DOLLAR__1905;
wire            n632____DOLLAR__1909;
wire            n633____DOLLAR__1913;
wire            n634____DOLLAR__1917;
wire            n635____DOLLAR__1921;
wire            n636____DOLLAR__1925;
wire            n637____DOLLAR__1929;
wire            n638____DOLLAR__1933;
wire            n639____DOLLAR__1937;
wire            n63____DOLLAR__321;
wire            n640____DOLLAR__1941;
wire            n641____DOLLAR__1945;
wire            n642____DOLLAR__1949;
wire            n643____DOLLAR__1953;
wire            n644____DOLLAR__1957;
wire            n645____DOLLAR__1961;
wire            n646____DOLLAR__1965;
wire            n647____DOLLAR__1969;
wire            n648____DOLLAR__1973;
wire            n649____DOLLAR__1977;
wire            n64____DOLLAR__325;
wire            n650____DOLLAR__1981;
wire            n651____DOLLAR__1985;
wire            n652____DOLLAR__1989;
wire            n653____DOLLAR__1993;
wire            n654____DOLLAR__1997;
wire            n655____DOLLAR__2001;
wire            n656____DOLLAR__2005;
wire            n657____DOLLAR__2009;
wire            n658____DOLLAR__2013;
wire            n659____DOLLAR__2017;
wire            n65____DOLLAR__329;
wire            n660____DOLLAR__2021;
wire            n661____DOLLAR__2025;
wire            n662____DOLLAR__2029;
wire            n663____DOLLAR__2033;
wire            n664____DOLLAR__2037;
wire            n665____DOLLAR__2041;
wire            n666____DOLLAR__2045;
wire            n667____DOLLAR__2049;
wire            n668____DOLLAR__2053;
wire            n669____DOLLAR__2057;
wire            n66____DOLLAR__333;
wire            n670____DOLLAR__2061;
wire            n671____DOLLAR__2065;
wire            n672____DOLLAR__2069;
wire            n673____DOLLAR__2073;
wire            n674____DOLLAR__2077;
wire            n675____DOLLAR__2081;
wire            n676____DOLLAR__2085;
wire            n677____DOLLAR__2089;
wire            n678____DOLLAR__2093;
wire            n679____DOLLAR__2097;
wire            n67____DOLLAR__337;
wire            n680____DOLLAR__2101;
wire            n681____DOLLAR__2105;
wire            n682____DOLLAR__2109;
wire            n683____DOLLAR__2113;
wire            n684____DOLLAR__2117;
wire            n685____DOLLAR__2121;
wire            n686____DOLLAR__2125;
wire            n687____DOLLAR__2129;
wire            n688____DOLLAR__2133;
wire            n689____DOLLAR__2137;
wire            n68____DOLLAR__341;
wire            n690____DOLLAR__2141;
wire            n691____DOLLAR__2143;
wire            n692____DOLLAR__2144;
wire            n693____DOLLAR__2145;
wire            n694____DOLLAR__2146;
wire            n695____DOLLAR__2147;
wire            n696____DOLLAR__2148;
wire            n697____DOLLAR__2149;
wire            n698____DOLLAR__2150;
wire            n699____DOLLAR__2151;
wire            n69____DOLLAR__345;
wire            n6____DOLLAR__93;
wire            n700____DOLLAR__2152;
wire            n701____DOLLAR__2153;
wire            n702____DOLLAR__2154;
wire            n703____DOLLAR__2155;
wire            n704____DOLLAR__2156;
wire            n705____DOLLAR__2157;
wire            n706____DOLLAR__2158;
wire            n707____DOLLAR__2159;
wire            n708____DOLLAR__2160;
wire            n709____DOLLAR__2161;
wire            n70____DOLLAR__349;
wire            n710____DOLLAR__2162;
wire            n711____DOLLAR__2163;
wire            n712____DOLLAR__2164;
wire            n713____DOLLAR__2165;
wire            n714____DOLLAR__2166;
wire            n715____DOLLAR__2167;
wire            n716____DOLLAR__2168;
wire            n717____DOLLAR__2169;
wire            n718____DOLLAR__2170;
wire            n719____DOLLAR__2171;
wire            n71____DOLLAR__353;
wire            n720____DOLLAR__2172;
wire            n721____DOLLAR__2173;
wire            n722____DOLLAR__2174;
wire            n723____DOLLAR__2175;
wire            n724____DOLLAR__2176;
wire            n725____DOLLAR__2177;
wire            n726____DOLLAR__2178;
wire            n727____DOLLAR__2179;
wire            n728____DOLLAR__2180;
wire            n729____DOLLAR__2181;
wire            n72____DOLLAR__357;
wire            n730____DOLLAR__2182;
wire            n731____DOLLAR__2183;
wire            n732____DOLLAR__2184;
wire            n733____DOLLAR__2185;
wire            n734____DOLLAR__2186;
wire            n735____DOLLAR__2187;
wire            n736____DOLLAR__2188;
wire            n737____DOLLAR__2189;
wire            n738____DOLLAR__2190;
wire            n739____DOLLAR__2191;
wire            n73____DOLLAR__361;
wire            n740____DOLLAR__2192;
wire            n741____DOLLAR__2193;
wire            n742____DOLLAR__2194;
wire            n743____DOLLAR__2195;
wire            n744____DOLLAR__2196;
wire            n745____DOLLAR__2197;
wire            n746____DOLLAR__2198;
wire            n747____DOLLAR__2199;
wire            n748____DOLLAR__2200;
wire            n749____DOLLAR__2201;
wire            n74____DOLLAR__365;
wire            n750____DOLLAR__2202;
wire            n751____DOLLAR__2203;
wire            n752____DOLLAR__2204;
wire            n753____DOLLAR__2205;
wire            n754____DOLLAR__2206;
wire            n755____DOLLAR__2207;
wire            n756____DOLLAR__2208;
wire            n757____DOLLAR__2209;
wire            n758____DOLLAR__2210;
wire            n759____DOLLAR__2211;
wire            n75____DOLLAR__369;
wire            n760____DOLLAR__2212;
wire            n761____DOLLAR__2213;
wire            n762____DOLLAR__2214;
wire            n763____DOLLAR__2215;
wire            n764____DOLLAR__2216;
wire            n765____DOLLAR__2217;
wire            n766____DOLLAR__2218;
wire            n767____DOLLAR__2219;
wire            n768____DOLLAR__2220;
wire            n769____DOLLAR__2221;
wire            n76____DOLLAR__373;
wire            n770____DOLLAR__2222;
wire            n771____DOLLAR__2223;
wire            n772____DOLLAR__2224;
wire            n773____DOLLAR__2225;
wire            n774____DOLLAR__2226;
wire            n775____DOLLAR__2227;
wire            n776____DOLLAR__2228;
wire            n777____DOLLAR__2229;
wire            n778____DOLLAR__2230;
wire            n779____DOLLAR__2231;
wire            n77____DOLLAR__377;
wire            n780____DOLLAR__2232;
wire            n781____DOLLAR__2233;
wire            n782____DOLLAR__2234;
wire            n783____DOLLAR__2235;
wire            n784____DOLLAR__2236;
wire            n785____DOLLAR__2237;
wire            n786____DOLLAR__2238;
wire            n787____DOLLAR__2239;
wire            n788____DOLLAR__2240;
wire            n789____DOLLAR__2241;
wire            n78____DOLLAR__381;
wire            n790____DOLLAR__2242;
wire            n791____DOLLAR__2243;
wire            n792____DOLLAR__2244;
wire            n793____DOLLAR__2245;
wire            n794____DOLLAR__2246;
wire            n795____DOLLAR__2247;
wire            n796____DOLLAR__2248;
wire            n797____DOLLAR__2249;
wire            n798____DOLLAR__2250;
wire            n799____DOLLAR__2251;
wire            n79____DOLLAR__385;
wire            n7____DOLLAR__97;
wire            n800____DOLLAR__2252;
wire            n801____DOLLAR__2253;
wire            n802____DOLLAR__2254;
wire            n803____DOLLAR__2255;
wire            n804____DOLLAR__2256;
wire            n805____DOLLAR__2257;
wire            n806____DOLLAR__2258;
wire            n807____DOLLAR__2259;
wire            n808____DOLLAR__2260;
wire            n809____DOLLAR__2261;
wire            n80____DOLLAR__389;
wire            n810____DOLLAR__2262;
wire            n811____DOLLAR__2263;
wire            n812____DOLLAR__2264;
wire            n813____DOLLAR__2265;
wire            n814____DOLLAR__2266;
wire            n815____DOLLAR__2267;
wire            n816____DOLLAR__2268;
wire            n817____DOLLAR__2269;
wire            n818____DOLLAR__2270;
wire            n819____DOLLAR__2271;
wire            n81____DOLLAR__393;
wire            n820____DOLLAR__2272;
wire            n821____DOLLAR__2273;
wire            n822____DOLLAR__2274;
wire            n823____DOLLAR__2275;
wire            n824____DOLLAR__2276;
wire            n825____DOLLAR__2277;
wire            n826____DOLLAR__2278;
wire            n827____DOLLAR__2279;
wire            n828____DOLLAR__2280;
wire            n829____DOLLAR__2281;
wire            n82____DOLLAR__397;
wire            n830____DOLLAR__2282;
wire            n831____DOLLAR__2283;
wire            n832____DOLLAR__2284;
wire            n833____DOLLAR__2285;
wire            n834____DOLLAR__2286;
wire            n835____DOLLAR__2287;
wire            n836____DOLLAR__2288;
wire            n837____DOLLAR__2289;
wire            n838____DOLLAR__2290;
wire            n839____DOLLAR__2291;
wire            n83____DOLLAR__401;
wire            n840____DOLLAR__2292;
wire            n841____DOLLAR__2293;
wire            n842____DOLLAR__2294;
wire            n843____DOLLAR__2295;
wire            n844____DOLLAR__2296;
wire            n845____DOLLAR__2297;
wire            n846____DOLLAR__2298;
wire            n847____DOLLAR__2299;
wire            n848____DOLLAR__2300;
wire            n849____DOLLAR__2301;
wire            n84____DOLLAR__405;
wire            n850____DOLLAR__2302;
wire            n851____DOLLAR__2303;
wire            n852____DOLLAR__2304;
wire            n853____DOLLAR__2305;
wire            n854____DOLLAR__2306;
wire            n855____DOLLAR__2307;
wire            n856____DOLLAR__2308;
wire            n857____DOLLAR__2309;
wire            n858____DOLLAR__2310;
wire            n859____DOLLAR__2311;
wire            n85____DOLLAR__409;
wire            n860____DOLLAR__2312;
wire            n861____DOLLAR__2313;
wire            n862____DOLLAR__2314;
wire            n863____DOLLAR__2315;
wire            n864____DOLLAR__2316;
wire            n865____DOLLAR__2317;
wire            n866____DOLLAR__2318;
wire            n867____DOLLAR__2319;
wire            n868____DOLLAR__2320;
wire            n869____DOLLAR__2321;
wire            n86____DOLLAR__413;
wire            n870____DOLLAR__2322;
wire            n871____DOLLAR__2323;
wire            n872____DOLLAR__2324;
wire            n873____DOLLAR__2325;
wire            n874____DOLLAR__2326;
wire            n875____DOLLAR__2327;
wire            n876____DOLLAR__2328;
wire            n877____DOLLAR__2329;
wire            n878____DOLLAR__2330;
wire            n879____DOLLAR__2331;
wire            n87____DOLLAR__417;
wire            n880____DOLLAR__2332;
wire            n881____DOLLAR__2333;
wire            n882____DOLLAR__2334;
wire            n883____DOLLAR__2335;
wire            n884____DOLLAR__2336;
wire            n885____DOLLAR__2337;
wire            n886____DOLLAR__2338;
wire            n887____DOLLAR__2339;
wire            n888____DOLLAR__2340;
wire            n889____DOLLAR__2341;
wire            n88____DOLLAR__421;
wire            n890____DOLLAR__2342;
wire            n891____DOLLAR__2343;
wire            n892____DOLLAR__2344;
wire            n893____DOLLAR__2345;
wire            n894____DOLLAR__2346;
wire            n895____DOLLAR__2347;
wire            n896____DOLLAR__2348;
wire            n897____DOLLAR__2349;
wire            n898____DOLLAR__2350;
wire            n899____DOLLAR__2351;
wire            n89____DOLLAR__425;
wire            n8____DOLLAR__101;
wire            n900____DOLLAR__2352;
wire            n901____DOLLAR__2353;
wire            n902____DOLLAR__2354;
wire            n903____DOLLAR__2355;
wire            n904____DOLLAR__2356;
wire            n905____DOLLAR__2357;
wire            n906____DOLLAR__2358;
wire            n907____DOLLAR__2359;
wire            n908____DOLLAR__2360;
wire            n909____DOLLAR__2361;
wire            n90____DOLLAR__429;
wire            n910____DOLLAR__2362;
wire            n911____DOLLAR__2363;
wire            n912____DOLLAR__2364;
wire            n913____DOLLAR__2365;
wire            n914____DOLLAR__2366;
wire            n915____DOLLAR__2367;
wire            n916____DOLLAR__2368;
wire      [1:0] n917____DOLLAR__2371;
wire      [4:0] n918____DOLLAR__2379;
wire      [7:0] n919____DOLLAR__2385;
wire            n91____DOLLAR__433;
wire            n920____DOLLAR__2389;
wire      [7:0] n921____DOLLAR__2391;
wire      [7:0] n922____DOLLAR__2392;
wire            n923____DOLLAR__2397;
wire            n924____DOLLAR__2401;
wire            n925____DOLLAR__2403;
wire      [3:0] n926____DOLLAR__177450;
wire            n927____DOLLAR__177531;
wire            n928____DOLLAR__177526;
wire            n929____DOLLAR__177521;
wire            n92____DOLLAR__437;
wire            n930____DOLLAR__177516;
wire            n931____DOLLAR__177511;
wire            n932____DOLLAR__177506;
wire            n933____DOLLAR__177501;
wire            n934____DOLLAR__177496;
wire            n935____DOLLAR__177491;
wire            n936____DOLLAR__177486;
wire            n937____DOLLAR__177481;
wire            n938____DOLLAR__177476;
wire            n939____DOLLAR__177471;
wire            n93____DOLLAR__441;
wire            n940____DOLLAR__177466;
wire            n941____DOLLAR__177461;
wire            n942____DOLLAR__177456;
wire      [7:0] n943____DOLLAR__177458;
wire      [7:0] n944____DOLLAR__177463;
wire      [7:0] n945____DOLLAR__177468;
wire      [7:0] n946____DOLLAR__177473;
wire      [7:0] n947____DOLLAR__177478;
wire      [7:0] n948____DOLLAR__177483;
wire      [7:0] n949____DOLLAR__177488;
wire            n94____DOLLAR__445;
wire      [7:0] n950____DOLLAR__177493;
wire      [7:0] n951____DOLLAR__177498;
wire      [7:0] n952____DOLLAR__177503;
wire      [7:0] n953____DOLLAR__177508;
wire      [7:0] n954____DOLLAR__177513;
wire      [7:0] n955____DOLLAR__177518;
wire      [7:0] n956____DOLLAR__177523;
wire      [7:0] n957____DOLLAR__177528;
wire      [7:0] n958____DOLLAR__177533;
wire      [7:0] n959____DOLLAR__2408;
wire            n95____DOLLAR__449;
wire      [3:0] n960____DOLLAR__177535;
wire            n961____DOLLAR__177616;
wire            n962____DOLLAR__177611;
wire            n963____DOLLAR__177606;
wire            n964____DOLLAR__177601;
wire            n965____DOLLAR__177596;
wire            n966____DOLLAR__177591;
wire            n967____DOLLAR__177586;
wire            n968____DOLLAR__177581;
wire            n969____DOLLAR__177576;
wire            n96____DOLLAR__453;
wire            n970____DOLLAR__177571;
wire            n971____DOLLAR__177566;
wire            n972____DOLLAR__177561;
wire            n973____DOLLAR__177556;
wire            n974____DOLLAR__177551;
wire            n975____DOLLAR__177546;
wire            n976____DOLLAR__177541;
wire      [7:0] n977____DOLLAR__177543;
wire      [7:0] n978____DOLLAR__177548;
wire      [7:0] n979____DOLLAR__177553;
wire            n97____DOLLAR__457;
wire      [7:0] n980____DOLLAR__177558;
wire      [7:0] n981____DOLLAR__177563;
wire      [7:0] n982____DOLLAR__177568;
wire      [7:0] n983____DOLLAR__177573;
wire      [7:0] n984____DOLLAR__177578;
wire      [7:0] n985____DOLLAR__177583;
wire      [7:0] n986____DOLLAR__177588;
wire      [7:0] n987____DOLLAR__177593;
wire      [7:0] n988____DOLLAR__177598;
wire      [7:0] n989____DOLLAR__177603;
wire            n98____DOLLAR__461;
wire      [7:0] n990____DOLLAR__177608;
wire      [7:0] n991____DOLLAR__177613;
wire      [7:0] n992____DOLLAR__177618;
wire     [15:0] n993____DOLLAR__2415;
wire            n994____DOLLAR__2421;
wire            n995____DOLLAR__2425;
wire            n996____DOLLAR__2427;
wire     [15:0] n997____DOLLAR__2430;
wire      [4:0] n998____DOLLAR__2431;
wire      [7:0] n999____DOLLAR__2439;
wire            n99____DOLLAR__465;
wire            n9____DOLLAR__105;
(* keep *) wire      [7:0] oc8051_IRAM_data_0_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_10_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_11_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_12_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_13_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_14_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_15_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_1_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_2_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_3_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_4_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_5_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_6_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_7_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_8_randinit;
(* keep *) wire      [7:0] oc8051_IRAM_data_9_randinit;
(* keep *) wire     [15:0] oc8051_ROM_addr_0_randinit;
(* keep *) wire     [15:0] oc8051_ROM_addr_1_randinit;
(* keep *) wire     [15:0] oc8051_ROM_addr_2_randinit;
wire      [7:0] oc8051_ROM_rdata_0;
wire      [7:0] oc8051_ROM_rdata_1;
wire      [7:0] oc8051_ROM_rdata_2;
wire            rst;
assign __ILA_oc8051_valid__ = 1'b1 ;
assign n0____DOLLAR__167758 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign __ILA_oc8051_decode_of_I__DOT__240__ = n0____DOLLAR__167758 ;
assign n2____DOLLAR__77 =  ( oc8051_ROM_rdata_0 ) == ( 8'd255 )  ;
assign n3____DOLLAR__81 =  ( oc8051_ROM_rdata_0 ) == ( 8'd254 )  ;
assign n4____DOLLAR__85 =  ( oc8051_ROM_rdata_0 ) == ( 8'd253 )  ;
assign n5____DOLLAR__89 =  ( oc8051_ROM_rdata_0 ) == ( 8'd252 )  ;
assign n6____DOLLAR__93 =  ( oc8051_ROM_rdata_0 ) == ( 8'd251 )  ;
assign n7____DOLLAR__97 =  ( oc8051_ROM_rdata_0 ) == ( 8'd250 )  ;
assign n8____DOLLAR__101 =  ( oc8051_ROM_rdata_0 ) == ( 8'd249 )  ;
assign n9____DOLLAR__105 =  ( oc8051_ROM_rdata_0 ) == ( 8'd248 )  ;
assign n10____DOLLAR__109 =  ( oc8051_ROM_rdata_0 ) == ( 8'd247 )  ;
assign n11____DOLLAR__113 =  ( oc8051_ROM_rdata_0 ) == ( 8'd246 )  ;
assign n12____DOLLAR__117 =  ( oc8051_ROM_rdata_0 ) == ( 8'd244 )  ;
assign n13____DOLLAR__121 =  ( oc8051_ROM_rdata_0 ) == ( 8'd243 )  ;
assign n14____DOLLAR__125 =  ( oc8051_ROM_rdata_0 ) == ( 8'd242 )  ;
assign n15____DOLLAR__129 =  ( oc8051_ROM_rdata_0 ) == ( 8'd241 )  ;
assign n16____DOLLAR__133 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign n17____DOLLAR__137 =  ( oc8051_ROM_rdata_0 ) == ( 8'd239 )  ;
assign n18____DOLLAR__141 =  ( oc8051_ROM_rdata_0 ) == ( 8'd238 )  ;
assign n19____DOLLAR__145 =  ( oc8051_ROM_rdata_0 ) == ( 8'd237 )  ;
assign n20____DOLLAR__149 =  ( oc8051_ROM_rdata_0 ) == ( 8'd236 )  ;
assign n21____DOLLAR__153 =  ( oc8051_ROM_rdata_0 ) == ( 8'd235 )  ;
assign n22____DOLLAR__157 =  ( oc8051_ROM_rdata_0 ) == ( 8'd234 )  ;
assign n23____DOLLAR__161 =  ( oc8051_ROM_rdata_0 ) == ( 8'd233 )  ;
assign n24____DOLLAR__165 =  ( oc8051_ROM_rdata_0 ) == ( 8'd232 )  ;
assign n25____DOLLAR__169 =  ( oc8051_ROM_rdata_0 ) == ( 8'd231 )  ;
assign n26____DOLLAR__173 =  ( oc8051_ROM_rdata_0 ) == ( 8'd230 )  ;
assign n27____DOLLAR__177 =  ( oc8051_ROM_rdata_0 ) == ( 8'd229 )  ;
assign n28____DOLLAR__181 =  ( oc8051_ROM_rdata_0 ) == ( 8'd228 )  ;
assign n29____DOLLAR__185 =  ( oc8051_ROM_rdata_0 ) == ( 8'd227 )  ;
assign n30____DOLLAR__189 =  ( oc8051_ROM_rdata_0 ) == ( 8'd226 )  ;
assign n31____DOLLAR__193 =  ( oc8051_ROM_rdata_0 ) == ( 8'd225 )  ;
assign n32____DOLLAR__197 =  ( oc8051_ROM_rdata_0 ) == ( 8'd224 )  ;
assign n33____DOLLAR__201 =  ( oc8051_ROM_rdata_0 ) == ( 8'd223 )  ;
assign n34____DOLLAR__205 =  ( oc8051_ROM_rdata_0 ) == ( 8'd222 )  ;
assign n35____DOLLAR__209 =  ( oc8051_ROM_rdata_0 ) == ( 8'd221 )  ;
assign n36____DOLLAR__213 =  ( oc8051_ROM_rdata_0 ) == ( 8'd220 )  ;
assign n37____DOLLAR__217 =  ( oc8051_ROM_rdata_0 ) == ( 8'd219 )  ;
assign n38____DOLLAR__221 =  ( oc8051_ROM_rdata_0 ) == ( 8'd218 )  ;
assign n39____DOLLAR__225 =  ( oc8051_ROM_rdata_0 ) == ( 8'd217 )  ;
assign n40____DOLLAR__229 =  ( oc8051_ROM_rdata_0 ) == ( 8'd216 )  ;
assign n41____DOLLAR__233 =  ( oc8051_ROM_rdata_0 ) == ( 8'd215 )  ;
assign n42____DOLLAR__237 =  ( oc8051_ROM_rdata_0 ) == ( 8'd214 )  ;
assign n43____DOLLAR__241 =  ( oc8051_ROM_rdata_0 ) == ( 8'd212 )  ;
assign n44____DOLLAR__245 =  ( oc8051_ROM_rdata_0 ) == ( 8'd211 )  ;
assign n45____DOLLAR__249 =  ( oc8051_ROM_rdata_0 ) == ( 8'd210 )  ;
assign n46____DOLLAR__253 =  ( oc8051_ROM_rdata_0 ) == ( 8'd209 )  ;
assign n47____DOLLAR__257 =  ( oc8051_ROM_rdata_0 ) == ( 8'd207 )  ;
assign n48____DOLLAR__261 =  ( oc8051_ROM_rdata_0 ) == ( 8'd206 )  ;
assign n49____DOLLAR__265 =  ( oc8051_ROM_rdata_0 ) == ( 8'd205 )  ;
assign n50____DOLLAR__269 =  ( oc8051_ROM_rdata_0 ) == ( 8'd204 )  ;
assign n51____DOLLAR__273 =  ( oc8051_ROM_rdata_0 ) == ( 8'd203 )  ;
assign n52____DOLLAR__277 =  ( oc8051_ROM_rdata_0 ) == ( 8'd202 )  ;
assign n53____DOLLAR__281 =  ( oc8051_ROM_rdata_0 ) == ( 8'd201 )  ;
assign n54____DOLLAR__285 =  ( oc8051_ROM_rdata_0 ) == ( 8'd200 )  ;
assign n55____DOLLAR__289 =  ( oc8051_ROM_rdata_0 ) == ( 8'd199 )  ;
assign n56____DOLLAR__293 =  ( oc8051_ROM_rdata_0 ) == ( 8'd198 )  ;
assign n57____DOLLAR__297 =  ( oc8051_ROM_rdata_0 ) == ( 8'd196 )  ;
assign n58____DOLLAR__301 =  ( oc8051_ROM_rdata_0 ) == ( 8'd195 )  ;
assign n59____DOLLAR__305 =  ( oc8051_ROM_rdata_0 ) == ( 8'd194 )  ;
assign n60____DOLLAR__309 =  ( oc8051_ROM_rdata_0 ) == ( 8'd193 )  ;
assign n61____DOLLAR__313 =  ( oc8051_ROM_rdata_0 ) == ( 8'd192 )  ;
assign n62____DOLLAR__317 =  ( oc8051_ROM_rdata_0 ) == ( 8'd191 )  ;
assign n63____DOLLAR__321 =  ( oc8051_ROM_rdata_0 ) == ( 8'd190 )  ;
assign n64____DOLLAR__325 =  ( oc8051_ROM_rdata_0 ) == ( 8'd189 )  ;
assign n65____DOLLAR__329 =  ( oc8051_ROM_rdata_0 ) == ( 8'd188 )  ;
assign n66____DOLLAR__333 =  ( oc8051_ROM_rdata_0 ) == ( 8'd187 )  ;
assign n67____DOLLAR__337 =  ( oc8051_ROM_rdata_0 ) == ( 8'd186 )  ;
assign n68____DOLLAR__341 =  ( oc8051_ROM_rdata_0 ) == ( 8'd185 )  ;
assign n69____DOLLAR__345 =  ( oc8051_ROM_rdata_0 ) == ( 8'd184 )  ;
assign n70____DOLLAR__349 =  ( oc8051_ROM_rdata_0 ) == ( 8'd183 )  ;
assign n71____DOLLAR__353 =  ( oc8051_ROM_rdata_0 ) == ( 8'd182 )  ;
assign n72____DOLLAR__357 =  ( oc8051_ROM_rdata_0 ) == ( 8'd181 )  ;
assign n73____DOLLAR__361 =  ( oc8051_ROM_rdata_0 ) == ( 8'd180 )  ;
assign n74____DOLLAR__365 =  ( oc8051_ROM_rdata_0 ) == ( 8'd179 )  ;
assign n75____DOLLAR__369 =  ( oc8051_ROM_rdata_0 ) == ( 8'd178 )  ;
assign n76____DOLLAR__373 =  ( oc8051_ROM_rdata_0 ) == ( 8'd177 )  ;
assign n77____DOLLAR__377 =  ( oc8051_ROM_rdata_0 ) == ( 8'd176 )  ;
assign n78____DOLLAR__381 =  ( oc8051_ROM_rdata_0 ) == ( 8'd175 )  ;
assign n79____DOLLAR__385 =  ( oc8051_ROM_rdata_0 ) == ( 8'd174 )  ;
assign n80____DOLLAR__389 =  ( oc8051_ROM_rdata_0 ) == ( 8'd173 )  ;
assign n81____DOLLAR__393 =  ( oc8051_ROM_rdata_0 ) == ( 8'd172 )  ;
assign n82____DOLLAR__397 =  ( oc8051_ROM_rdata_0 ) == ( 8'd171 )  ;
assign n83____DOLLAR__401 =  ( oc8051_ROM_rdata_0 ) == ( 8'd170 )  ;
assign n84____DOLLAR__405 =  ( oc8051_ROM_rdata_0 ) == ( 8'd169 )  ;
assign n85____DOLLAR__409 =  ( oc8051_ROM_rdata_0 ) == ( 8'd168 )  ;
assign n86____DOLLAR__413 =  ( oc8051_ROM_rdata_0 ) == ( 8'd167 )  ;
assign n87____DOLLAR__417 =  ( oc8051_ROM_rdata_0 ) == ( 8'd166 )  ;
assign n88____DOLLAR__421 =  ( oc8051_ROM_rdata_0 ) == ( 8'd165 )  ;
assign n89____DOLLAR__425 =  ( oc8051_ROM_rdata_0 ) == ( 8'd164 )  ;
assign n90____DOLLAR__429 =  ( oc8051_ROM_rdata_0 ) == ( 8'd162 )  ;
assign n91____DOLLAR__433 =  ( oc8051_ROM_rdata_0 ) == ( 8'd161 )  ;
assign n92____DOLLAR__437 =  ( oc8051_ROM_rdata_0 ) == ( 8'd160 )  ;
assign n93____DOLLAR__441 =  ( oc8051_ROM_rdata_0 ) == ( 8'd159 )  ;
assign n94____DOLLAR__445 =  ( oc8051_ROM_rdata_0 ) == ( 8'd158 )  ;
assign n95____DOLLAR__449 =  ( oc8051_ROM_rdata_0 ) == ( 8'd157 )  ;
assign n96____DOLLAR__453 =  ( oc8051_ROM_rdata_0 ) == ( 8'd156 )  ;
assign n97____DOLLAR__457 =  ( oc8051_ROM_rdata_0 ) == ( 8'd155 )  ;
assign n98____DOLLAR__461 =  ( oc8051_ROM_rdata_0 ) == ( 8'd154 )  ;
assign n99____DOLLAR__465 =  ( oc8051_ROM_rdata_0 ) == ( 8'd153 )  ;
assign n100____DOLLAR__469 =  ( oc8051_ROM_rdata_0 ) == ( 8'd152 )  ;
assign n101____DOLLAR__473 =  ( oc8051_ROM_rdata_0 ) == ( 8'd151 )  ;
assign n102____DOLLAR__477 =  ( oc8051_ROM_rdata_0 ) == ( 8'd150 )  ;
assign n103____DOLLAR__481 =  ( oc8051_ROM_rdata_0 ) == ( 8'd149 )  ;
assign n104____DOLLAR__485 =  ( oc8051_ROM_rdata_0 ) == ( 8'd148 )  ;
assign n105____DOLLAR__489 =  ( oc8051_ROM_rdata_0 ) == ( 8'd147 )  ;
assign n106____DOLLAR__493 =  ( oc8051_ROM_rdata_0 ) == ( 8'd146 )  ;
assign n107____DOLLAR__497 =  ( oc8051_ROM_rdata_0 ) == ( 8'd145 )  ;
assign n108____DOLLAR__501 =  ( oc8051_ROM_rdata_0 ) == ( 8'd132 )  ;
assign n109____DOLLAR__505 =  ( oc8051_ROM_rdata_0 ) == ( 8'd131 )  ;
assign n110____DOLLAR__509 =  ( oc8051_ROM_rdata_0 ) == ( 8'd130 )  ;
assign n111____DOLLAR__513 =  ( oc8051_ROM_rdata_0 ) == ( 8'd129 )  ;
assign n112____DOLLAR__517 =  ( oc8051_ROM_rdata_0 ) == ( 8'd128 )  ;
assign n113____DOLLAR__521 =  ( oc8051_ROM_rdata_0 ) == ( 8'd127 )  ;
assign n114____DOLLAR__525 =  ( oc8051_ROM_rdata_0 ) == ( 8'd126 )  ;
assign n115____DOLLAR__529 =  ( oc8051_ROM_rdata_0 ) == ( 8'd125 )  ;
assign n116____DOLLAR__533 =  ( oc8051_ROM_rdata_0 ) == ( 8'd124 )  ;
assign n117____DOLLAR__537 =  ( oc8051_ROM_rdata_0 ) == ( 8'd123 )  ;
assign n118____DOLLAR__541 =  ( oc8051_ROM_rdata_0 ) == ( 8'd122 )  ;
assign n119____DOLLAR__545 =  ( oc8051_ROM_rdata_0 ) == ( 8'd121 )  ;
assign n120____DOLLAR__549 =  ( oc8051_ROM_rdata_0 ) == ( 8'd120 )  ;
assign n121____DOLLAR__553 =  ( oc8051_ROM_rdata_0 ) == ( 8'd119 )  ;
assign n122____DOLLAR__557 =  ( oc8051_ROM_rdata_0 ) == ( 8'd118 )  ;
assign n123____DOLLAR__561 =  ( oc8051_ROM_rdata_0 ) == ( 8'd116 )  ;
assign n124____DOLLAR__565 =  ( oc8051_ROM_rdata_0 ) == ( 8'd115 )  ;
assign n125____DOLLAR__569 =  ( oc8051_ROM_rdata_0 ) == ( 8'd114 )  ;
assign n126____DOLLAR__573 =  ( oc8051_ROM_rdata_0 ) == ( 8'd113 )  ;
assign n127____DOLLAR__577 =  ( oc8051_ROM_rdata_0 ) == ( 8'd112 )  ;
assign n128____DOLLAR__581 =  ( oc8051_ROM_rdata_0 ) == ( 8'd111 )  ;
assign n129____DOLLAR__585 =  ( oc8051_ROM_rdata_0 ) == ( 8'd110 )  ;
assign n130____DOLLAR__589 =  ( oc8051_ROM_rdata_0 ) == ( 8'd109 )  ;
assign n131____DOLLAR__593 =  ( oc8051_ROM_rdata_0 ) == ( 8'd108 )  ;
assign n132____DOLLAR__597 =  ( oc8051_ROM_rdata_0 ) == ( 8'd107 )  ;
assign n133____DOLLAR__601 =  ( oc8051_ROM_rdata_0 ) == ( 8'd106 )  ;
assign n134____DOLLAR__605 =  ( oc8051_ROM_rdata_0 ) == ( 8'd105 )  ;
assign n135____DOLLAR__609 =  ( oc8051_ROM_rdata_0 ) == ( 8'd104 )  ;
assign n136____DOLLAR__613 =  ( oc8051_ROM_rdata_0 ) == ( 8'd103 )  ;
assign n137____DOLLAR__617 =  ( oc8051_ROM_rdata_0 ) == ( 8'd102 )  ;
assign n138____DOLLAR__621 =  ( oc8051_ROM_rdata_0 ) == ( 8'd101 )  ;
assign n139____DOLLAR__625 =  ( oc8051_ROM_rdata_0 ) == ( 8'd100 )  ;
assign n140____DOLLAR__629 =  ( oc8051_ROM_rdata_0 ) == ( 8'd97 )  ;
assign n141____DOLLAR__633 =  ( oc8051_ROM_rdata_0 ) == ( 8'd96 )  ;
assign n142____DOLLAR__637 =  ( oc8051_ROM_rdata_0 ) == ( 8'd95 )  ;
assign n143____DOLLAR__641 =  ( oc8051_ROM_rdata_0 ) == ( 8'd94 )  ;
assign n144____DOLLAR__645 =  ( oc8051_ROM_rdata_0 ) == ( 8'd93 )  ;
assign n145____DOLLAR__649 =  ( oc8051_ROM_rdata_0 ) == ( 8'd92 )  ;
assign n146____DOLLAR__653 =  ( oc8051_ROM_rdata_0 ) == ( 8'd91 )  ;
assign n147____DOLLAR__657 =  ( oc8051_ROM_rdata_0 ) == ( 8'd90 )  ;
assign n148____DOLLAR__661 =  ( oc8051_ROM_rdata_0 ) == ( 8'd89 )  ;
assign n149____DOLLAR__665 =  ( oc8051_ROM_rdata_0 ) == ( 8'd88 )  ;
assign n150____DOLLAR__669 =  ( oc8051_ROM_rdata_0 ) == ( 8'd87 )  ;
assign n151____DOLLAR__673 =  ( oc8051_ROM_rdata_0 ) == ( 8'd86 )  ;
assign n152____DOLLAR__677 =  ( oc8051_ROM_rdata_0 ) == ( 8'd85 )  ;
assign n153____DOLLAR__681 =  ( oc8051_ROM_rdata_0 ) == ( 8'd84 )  ;
assign n154____DOLLAR__685 =  ( oc8051_ROM_rdata_0 ) == ( 8'd81 )  ;
assign n155____DOLLAR__689 =  ( oc8051_ROM_rdata_0 ) == ( 8'd80 )  ;
assign n156____DOLLAR__693 =  ( oc8051_ROM_rdata_0 ) == ( 8'd79 )  ;
assign n157____DOLLAR__697 =  ( oc8051_ROM_rdata_0 ) == ( 8'd78 )  ;
assign n158____DOLLAR__701 =  ( oc8051_ROM_rdata_0 ) == ( 8'd77 )  ;
assign n159____DOLLAR__705 =  ( oc8051_ROM_rdata_0 ) == ( 8'd76 )  ;
assign n160____DOLLAR__709 =  ( oc8051_ROM_rdata_0 ) == ( 8'd75 )  ;
assign n161____DOLLAR__713 =  ( oc8051_ROM_rdata_0 ) == ( 8'd74 )  ;
assign n162____DOLLAR__717 =  ( oc8051_ROM_rdata_0 ) == ( 8'd73 )  ;
assign n163____DOLLAR__721 =  ( oc8051_ROM_rdata_0 ) == ( 8'd72 )  ;
assign n164____DOLLAR__725 =  ( oc8051_ROM_rdata_0 ) == ( 8'd71 )  ;
assign n165____DOLLAR__729 =  ( oc8051_ROM_rdata_0 ) == ( 8'd70 )  ;
assign n166____DOLLAR__733 =  ( oc8051_ROM_rdata_0 ) == ( 8'd69 )  ;
assign n167____DOLLAR__737 =  ( oc8051_ROM_rdata_0 ) == ( 8'd68 )  ;
assign n168____DOLLAR__741 =  ( oc8051_ROM_rdata_0 ) == ( 8'd65 )  ;
assign n169____DOLLAR__745 =  ( oc8051_ROM_rdata_0 ) == ( 8'd64 )  ;
assign n170____DOLLAR__749 =  ( oc8051_ROM_rdata_0 ) == ( 8'd63 )  ;
assign n171____DOLLAR__753 =  ( oc8051_ROM_rdata_0 ) == ( 8'd62 )  ;
assign n172____DOLLAR__757 =  ( oc8051_ROM_rdata_0 ) == ( 8'd61 )  ;
assign n173____DOLLAR__761 =  ( oc8051_ROM_rdata_0 ) == ( 8'd60 )  ;
assign n174____DOLLAR__765 =  ( oc8051_ROM_rdata_0 ) == ( 8'd59 )  ;
assign n175____DOLLAR__769 =  ( oc8051_ROM_rdata_0 ) == ( 8'd58 )  ;
assign n176____DOLLAR__773 =  ( oc8051_ROM_rdata_0 ) == ( 8'd57 )  ;
assign n177____DOLLAR__777 =  ( oc8051_ROM_rdata_0 ) == ( 8'd56 )  ;
assign n178____DOLLAR__781 =  ( oc8051_ROM_rdata_0 ) == ( 8'd55 )  ;
assign n179____DOLLAR__785 =  ( oc8051_ROM_rdata_0 ) == ( 8'd54 )  ;
assign n180____DOLLAR__789 =  ( oc8051_ROM_rdata_0 ) == ( 8'd53 )  ;
assign n181____DOLLAR__793 =  ( oc8051_ROM_rdata_0 ) == ( 8'd52 )  ;
assign n182____DOLLAR__797 =  ( oc8051_ROM_rdata_0 ) == ( 8'd51 )  ;
assign n183____DOLLAR__801 =  ( oc8051_ROM_rdata_0 ) == ( 8'd50 )  ;
assign n184____DOLLAR__805 =  ( oc8051_ROM_rdata_0 ) == ( 8'd49 )  ;
assign n185____DOLLAR__809 =  ( oc8051_ROM_rdata_0 ) == ( 8'd48 )  ;
assign n186____DOLLAR__813 =  ( oc8051_ROM_rdata_0 ) == ( 8'd47 )  ;
assign n187____DOLLAR__817 =  ( oc8051_ROM_rdata_0 ) == ( 8'd46 )  ;
assign n188____DOLLAR__821 =  ( oc8051_ROM_rdata_0 ) == ( 8'd45 )  ;
assign n189____DOLLAR__825 =  ( oc8051_ROM_rdata_0 ) == ( 8'd44 )  ;
assign n190____DOLLAR__829 =  ( oc8051_ROM_rdata_0 ) == ( 8'd43 )  ;
assign n191____DOLLAR__833 =  ( oc8051_ROM_rdata_0 ) == ( 8'd42 )  ;
assign n192____DOLLAR__837 =  ( oc8051_ROM_rdata_0 ) == ( 8'd41 )  ;
assign n193____DOLLAR__841 =  ( oc8051_ROM_rdata_0 ) == ( 8'd40 )  ;
assign n194____DOLLAR__845 =  ( oc8051_ROM_rdata_0 ) == ( 8'd39 )  ;
assign n195____DOLLAR__849 =  ( oc8051_ROM_rdata_0 ) == ( 8'd38 )  ;
assign n196____DOLLAR__853 =  ( oc8051_ROM_rdata_0 ) == ( 8'd37 )  ;
assign n197____DOLLAR__857 =  ( oc8051_ROM_rdata_0 ) == ( 8'd36 )  ;
assign n198____DOLLAR__861 =  ( oc8051_ROM_rdata_0 ) == ( 8'd35 )  ;
assign n199____DOLLAR__865 =  ( oc8051_ROM_rdata_0 ) == ( 8'd34 )  ;
assign n200____DOLLAR__869 =  ( oc8051_ROM_rdata_0 ) == ( 8'd33 )  ;
assign n201____DOLLAR__873 =  ( oc8051_ROM_rdata_0 ) == ( 8'd32 )  ;
assign n202____DOLLAR__877 =  ( oc8051_ROM_rdata_0 ) == ( 8'd31 )  ;
assign n203____DOLLAR__881 =  ( oc8051_ROM_rdata_0 ) == ( 8'd30 )  ;
assign n204____DOLLAR__885 =  ( oc8051_ROM_rdata_0 ) == ( 8'd29 )  ;
assign n205____DOLLAR__889 =  ( oc8051_ROM_rdata_0 ) == ( 8'd28 )  ;
assign n206____DOLLAR__893 =  ( oc8051_ROM_rdata_0 ) == ( 8'd27 )  ;
assign n207____DOLLAR__897 =  ( oc8051_ROM_rdata_0 ) == ( 8'd26 )  ;
assign n208____DOLLAR__901 =  ( oc8051_ROM_rdata_0 ) == ( 8'd25 )  ;
assign n209____DOLLAR__905 =  ( oc8051_ROM_rdata_0 ) == ( 8'd24 )  ;
assign n210____DOLLAR__909 =  ( oc8051_ROM_rdata_0 ) == ( 8'd23 )  ;
assign n211____DOLLAR__913 =  ( oc8051_ROM_rdata_0 ) == ( 8'd22 )  ;
assign n212____DOLLAR__917 =  ( oc8051_ROM_rdata_0 ) == ( 8'd20 )  ;
assign n213____DOLLAR__921 =  ( oc8051_ROM_rdata_0 ) == ( 8'd19 )  ;
assign n214____DOLLAR__925 =  ( oc8051_ROM_rdata_0 ) == ( 8'd18 )  ;
assign n215____DOLLAR__929 =  ( oc8051_ROM_rdata_0 ) == ( 8'd17 )  ;
assign n216____DOLLAR__933 =  ( oc8051_ROM_rdata_0 ) == ( 8'd16 )  ;
assign n217____DOLLAR__937 =  ( oc8051_ROM_rdata_0 ) == ( 8'd15 )  ;
assign n218____DOLLAR__941 =  ( oc8051_ROM_rdata_0 ) == ( 8'd14 )  ;
assign n219____DOLLAR__945 =  ( oc8051_ROM_rdata_0 ) == ( 8'd13 )  ;
assign n220____DOLLAR__949 =  ( oc8051_ROM_rdata_0 ) == ( 8'd12 )  ;
assign n221____DOLLAR__953 =  ( oc8051_ROM_rdata_0 ) == ( 8'd11 )  ;
assign n222____DOLLAR__957 =  ( oc8051_ROM_rdata_0 ) == ( 8'd10 )  ;
assign n223____DOLLAR__961 =  ( oc8051_ROM_rdata_0 ) == ( 8'd9 )  ;
assign n224____DOLLAR__965 =  ( oc8051_ROM_rdata_0 ) == ( 8'd8 )  ;
assign n225____DOLLAR__969 =  ( oc8051_ROM_rdata_0 ) == ( 8'd7 )  ;
assign n226____DOLLAR__973 =  ( oc8051_ROM_rdata_0 ) == ( 8'd6 )  ;
assign n227____DOLLAR__977 =  ( oc8051_ROM_rdata_0 ) == ( 8'd4 )  ;
assign n228____DOLLAR__981 =  ( oc8051_ROM_rdata_0 ) == ( 8'd3 )  ;
assign n229____DOLLAR__985 =  ( oc8051_ROM_rdata_0 ) == ( 8'd2 )  ;
assign n230____DOLLAR__989 =  ( oc8051_ROM_rdata_0 ) == ( 8'd1 )  ;
assign n231____DOLLAR__993 =  ( oc8051_ROM_rdata_0 ) == ( 8'd0 )  ;
assign n232____DOLLAR__995 =  ( n230____DOLLAR__989 ) | ( n231____DOLLAR__993 )  ;
assign n233____DOLLAR__996 =  ( n229____DOLLAR__985 ) | ( n232____DOLLAR__995 )  ;
assign n234____DOLLAR__997 =  ( n228____DOLLAR__981 ) | ( n233____DOLLAR__996 )  ;
assign n235____DOLLAR__998 =  ( n227____DOLLAR__977 ) | ( n234____DOLLAR__997 )  ;
assign n236____DOLLAR__999 =  ( n226____DOLLAR__973 ) | ( n235____DOLLAR__998 )  ;
assign n237____DOLLAR__1000 =  ( n225____DOLLAR__969 ) | ( n236____DOLLAR__999 )  ;
assign n238____DOLLAR__1001 =  ( n224____DOLLAR__965 ) | ( n237____DOLLAR__1000 )  ;
assign n239____DOLLAR__1002 =  ( n223____DOLLAR__961 ) | ( n238____DOLLAR__1001 )  ;
assign n240____DOLLAR__1003 =  ( n222____DOLLAR__957 ) | ( n239____DOLLAR__1002 )  ;
assign n241____DOLLAR__1004 =  ( n221____DOLLAR__953 ) | ( n240____DOLLAR__1003 )  ;
assign n242____DOLLAR__1005 =  ( n220____DOLLAR__949 ) | ( n241____DOLLAR__1004 )  ;
assign n243____DOLLAR__1006 =  ( n219____DOLLAR__945 ) | ( n242____DOLLAR__1005 )  ;
assign n244____DOLLAR__1007 =  ( n218____DOLLAR__941 ) | ( n243____DOLLAR__1006 )  ;
assign n245____DOLLAR__1008 =  ( n217____DOLLAR__937 ) | ( n244____DOLLAR__1007 )  ;
assign n246____DOLLAR__1009 =  ( n216____DOLLAR__933 ) | ( n245____DOLLAR__1008 )  ;
assign n247____DOLLAR__1010 =  ( n215____DOLLAR__929 ) | ( n246____DOLLAR__1009 )  ;
assign n248____DOLLAR__1011 =  ( n214____DOLLAR__925 ) | ( n247____DOLLAR__1010 )  ;
assign n249____DOLLAR__1012 =  ( n213____DOLLAR__921 ) | ( n248____DOLLAR__1011 )  ;
assign n250____DOLLAR__1013 =  ( n212____DOLLAR__917 ) | ( n249____DOLLAR__1012 )  ;
assign n251____DOLLAR__1014 =  ( n211____DOLLAR__913 ) | ( n250____DOLLAR__1013 )  ;
assign n252____DOLLAR__1015 =  ( n210____DOLLAR__909 ) | ( n251____DOLLAR__1014 )  ;
assign n253____DOLLAR__1016 =  ( n209____DOLLAR__905 ) | ( n252____DOLLAR__1015 )  ;
assign n254____DOLLAR__1017 =  ( n208____DOLLAR__901 ) | ( n253____DOLLAR__1016 )  ;
assign n255____DOLLAR__1018 =  ( n207____DOLLAR__897 ) | ( n254____DOLLAR__1017 )  ;
assign n256____DOLLAR__1019 =  ( n206____DOLLAR__893 ) | ( n255____DOLLAR__1018 )  ;
assign n257____DOLLAR__1020 =  ( n205____DOLLAR__889 ) | ( n256____DOLLAR__1019 )  ;
assign n258____DOLLAR__1021 =  ( n204____DOLLAR__885 ) | ( n257____DOLLAR__1020 )  ;
assign n259____DOLLAR__1022 =  ( n203____DOLLAR__881 ) | ( n258____DOLLAR__1021 )  ;
assign n260____DOLLAR__1023 =  ( n202____DOLLAR__877 ) | ( n259____DOLLAR__1022 )  ;
assign n261____DOLLAR__1024 =  ( n201____DOLLAR__873 ) | ( n260____DOLLAR__1023 )  ;
assign n262____DOLLAR__1025 =  ( n200____DOLLAR__869 ) | ( n261____DOLLAR__1024 )  ;
assign n263____DOLLAR__1026 =  ( n199____DOLLAR__865 ) | ( n262____DOLLAR__1025 )  ;
assign n264____DOLLAR__1027 =  ( n198____DOLLAR__861 ) | ( n263____DOLLAR__1026 )  ;
assign n265____DOLLAR__1028 =  ( n197____DOLLAR__857 ) | ( n264____DOLLAR__1027 )  ;
assign n266____DOLLAR__1029 =  ( n196____DOLLAR__853 ) | ( n265____DOLLAR__1028 )  ;
assign n267____DOLLAR__1030 =  ( n195____DOLLAR__849 ) | ( n266____DOLLAR__1029 )  ;
assign n268____DOLLAR__1031 =  ( n194____DOLLAR__845 ) | ( n267____DOLLAR__1030 )  ;
assign n269____DOLLAR__1032 =  ( n193____DOLLAR__841 ) | ( n268____DOLLAR__1031 )  ;
assign n270____DOLLAR__1033 =  ( n192____DOLLAR__837 ) | ( n269____DOLLAR__1032 )  ;
assign n271____DOLLAR__1034 =  ( n191____DOLLAR__833 ) | ( n270____DOLLAR__1033 )  ;
assign n272____DOLLAR__1035 =  ( n190____DOLLAR__829 ) | ( n271____DOLLAR__1034 )  ;
assign n273____DOLLAR__1036 =  ( n189____DOLLAR__825 ) | ( n272____DOLLAR__1035 )  ;
assign n274____DOLLAR__1037 =  ( n188____DOLLAR__821 ) | ( n273____DOLLAR__1036 )  ;
assign n275____DOLLAR__1038 =  ( n187____DOLLAR__817 ) | ( n274____DOLLAR__1037 )  ;
assign n276____DOLLAR__1039 =  ( n186____DOLLAR__813 ) | ( n275____DOLLAR__1038 )  ;
assign n277____DOLLAR__1040 =  ( n185____DOLLAR__809 ) | ( n276____DOLLAR__1039 )  ;
assign n278____DOLLAR__1041 =  ( n184____DOLLAR__805 ) | ( n277____DOLLAR__1040 )  ;
assign n279____DOLLAR__1042 =  ( n183____DOLLAR__801 ) | ( n278____DOLLAR__1041 )  ;
assign n280____DOLLAR__1043 =  ( n182____DOLLAR__797 ) | ( n279____DOLLAR__1042 )  ;
assign n281____DOLLAR__1044 =  ( n181____DOLLAR__793 ) | ( n280____DOLLAR__1043 )  ;
assign n282____DOLLAR__1045 =  ( n180____DOLLAR__789 ) | ( n281____DOLLAR__1044 )  ;
assign n283____DOLLAR__1046 =  ( n179____DOLLAR__785 ) | ( n282____DOLLAR__1045 )  ;
assign n284____DOLLAR__1047 =  ( n178____DOLLAR__781 ) | ( n283____DOLLAR__1046 )  ;
assign n285____DOLLAR__1048 =  ( n177____DOLLAR__777 ) | ( n284____DOLLAR__1047 )  ;
assign n286____DOLLAR__1049 =  ( n176____DOLLAR__773 ) | ( n285____DOLLAR__1048 )  ;
assign n287____DOLLAR__1050 =  ( n175____DOLLAR__769 ) | ( n286____DOLLAR__1049 )  ;
assign n288____DOLLAR__1051 =  ( n174____DOLLAR__765 ) | ( n287____DOLLAR__1050 )  ;
assign n289____DOLLAR__1052 =  ( n173____DOLLAR__761 ) | ( n288____DOLLAR__1051 )  ;
assign n290____DOLLAR__1053 =  ( n172____DOLLAR__757 ) | ( n289____DOLLAR__1052 )  ;
assign n291____DOLLAR__1054 =  ( n171____DOLLAR__753 ) | ( n290____DOLLAR__1053 )  ;
assign n292____DOLLAR__1055 =  ( n170____DOLLAR__749 ) | ( n291____DOLLAR__1054 )  ;
assign n293____DOLLAR__1056 =  ( n169____DOLLAR__745 ) | ( n292____DOLLAR__1055 )  ;
assign n294____DOLLAR__1057 =  ( n168____DOLLAR__741 ) | ( n293____DOLLAR__1056 )  ;
assign n295____DOLLAR__1058 =  ( n167____DOLLAR__737 ) | ( n294____DOLLAR__1057 )  ;
assign n296____DOLLAR__1059 =  ( n166____DOLLAR__733 ) | ( n295____DOLLAR__1058 )  ;
assign n297____DOLLAR__1060 =  ( n165____DOLLAR__729 ) | ( n296____DOLLAR__1059 )  ;
assign n298____DOLLAR__1061 =  ( n164____DOLLAR__725 ) | ( n297____DOLLAR__1060 )  ;
assign n299____DOLLAR__1062 =  ( n163____DOLLAR__721 ) | ( n298____DOLLAR__1061 )  ;
assign n300____DOLLAR__1063 =  ( n162____DOLLAR__717 ) | ( n299____DOLLAR__1062 )  ;
assign n301____DOLLAR__1064 =  ( n161____DOLLAR__713 ) | ( n300____DOLLAR__1063 )  ;
assign n302____DOLLAR__1065 =  ( n160____DOLLAR__709 ) | ( n301____DOLLAR__1064 )  ;
assign n303____DOLLAR__1066 =  ( n159____DOLLAR__705 ) | ( n302____DOLLAR__1065 )  ;
assign n304____DOLLAR__1067 =  ( n158____DOLLAR__701 ) | ( n303____DOLLAR__1066 )  ;
assign n305____DOLLAR__1068 =  ( n157____DOLLAR__697 ) | ( n304____DOLLAR__1067 )  ;
assign n306____DOLLAR__1069 =  ( n156____DOLLAR__693 ) | ( n305____DOLLAR__1068 )  ;
assign n307____DOLLAR__1070 =  ( n155____DOLLAR__689 ) | ( n306____DOLLAR__1069 )  ;
assign n308____DOLLAR__1071 =  ( n154____DOLLAR__685 ) | ( n307____DOLLAR__1070 )  ;
assign n309____DOLLAR__1072 =  ( n153____DOLLAR__681 ) | ( n308____DOLLAR__1071 )  ;
assign n310____DOLLAR__1073 =  ( n152____DOLLAR__677 ) | ( n309____DOLLAR__1072 )  ;
assign n311____DOLLAR__1074 =  ( n151____DOLLAR__673 ) | ( n310____DOLLAR__1073 )  ;
assign n312____DOLLAR__1075 =  ( n150____DOLLAR__669 ) | ( n311____DOLLAR__1074 )  ;
assign n313____DOLLAR__1076 =  ( n149____DOLLAR__665 ) | ( n312____DOLLAR__1075 )  ;
assign n314____DOLLAR__1077 =  ( n148____DOLLAR__661 ) | ( n313____DOLLAR__1076 )  ;
assign n315____DOLLAR__1078 =  ( n147____DOLLAR__657 ) | ( n314____DOLLAR__1077 )  ;
assign n316____DOLLAR__1079 =  ( n146____DOLLAR__653 ) | ( n315____DOLLAR__1078 )  ;
assign n317____DOLLAR__1080 =  ( n145____DOLLAR__649 ) | ( n316____DOLLAR__1079 )  ;
assign n318____DOLLAR__1081 =  ( n144____DOLLAR__645 ) | ( n317____DOLLAR__1080 )  ;
assign n319____DOLLAR__1082 =  ( n143____DOLLAR__641 ) | ( n318____DOLLAR__1081 )  ;
assign n320____DOLLAR__1083 =  ( n142____DOLLAR__637 ) | ( n319____DOLLAR__1082 )  ;
assign n321____DOLLAR__1084 =  ( n141____DOLLAR__633 ) | ( n320____DOLLAR__1083 )  ;
assign n322____DOLLAR__1085 =  ( n140____DOLLAR__629 ) | ( n321____DOLLAR__1084 )  ;
assign n323____DOLLAR__1086 =  ( n139____DOLLAR__625 ) | ( n322____DOLLAR__1085 )  ;
assign n324____DOLLAR__1087 =  ( n138____DOLLAR__621 ) | ( n323____DOLLAR__1086 )  ;
assign n325____DOLLAR__1088 =  ( n137____DOLLAR__617 ) | ( n324____DOLLAR__1087 )  ;
assign n326____DOLLAR__1089 =  ( n136____DOLLAR__613 ) | ( n325____DOLLAR__1088 )  ;
assign n327____DOLLAR__1090 =  ( n135____DOLLAR__609 ) | ( n326____DOLLAR__1089 )  ;
assign n328____DOLLAR__1091 =  ( n134____DOLLAR__605 ) | ( n327____DOLLAR__1090 )  ;
assign n329____DOLLAR__1092 =  ( n133____DOLLAR__601 ) | ( n328____DOLLAR__1091 )  ;
assign n330____DOLLAR__1093 =  ( n132____DOLLAR__597 ) | ( n329____DOLLAR__1092 )  ;
assign n331____DOLLAR__1094 =  ( n131____DOLLAR__593 ) | ( n330____DOLLAR__1093 )  ;
assign n332____DOLLAR__1095 =  ( n130____DOLLAR__589 ) | ( n331____DOLLAR__1094 )  ;
assign n333____DOLLAR__1096 =  ( n129____DOLLAR__585 ) | ( n332____DOLLAR__1095 )  ;
assign n334____DOLLAR__1097 =  ( n128____DOLLAR__581 ) | ( n333____DOLLAR__1096 )  ;
assign n335____DOLLAR__1098 =  ( n127____DOLLAR__577 ) | ( n334____DOLLAR__1097 )  ;
assign n336____DOLLAR__1099 =  ( n126____DOLLAR__573 ) | ( n335____DOLLAR__1098 )  ;
assign n337____DOLLAR__1100 =  ( n125____DOLLAR__569 ) | ( n336____DOLLAR__1099 )  ;
assign n338____DOLLAR__1101 =  ( n124____DOLLAR__565 ) | ( n337____DOLLAR__1100 )  ;
assign n339____DOLLAR__1102 =  ( n123____DOLLAR__561 ) | ( n338____DOLLAR__1101 )  ;
assign n340____DOLLAR__1103 =  ( n122____DOLLAR__557 ) | ( n339____DOLLAR__1102 )  ;
assign n341____DOLLAR__1104 =  ( n121____DOLLAR__553 ) | ( n340____DOLLAR__1103 )  ;
assign n342____DOLLAR__1105 =  ( n120____DOLLAR__549 ) | ( n341____DOLLAR__1104 )  ;
assign n343____DOLLAR__1106 =  ( n119____DOLLAR__545 ) | ( n342____DOLLAR__1105 )  ;
assign n344____DOLLAR__1107 =  ( n118____DOLLAR__541 ) | ( n343____DOLLAR__1106 )  ;
assign n345____DOLLAR__1108 =  ( n117____DOLLAR__537 ) | ( n344____DOLLAR__1107 )  ;
assign n346____DOLLAR__1109 =  ( n116____DOLLAR__533 ) | ( n345____DOLLAR__1108 )  ;
assign n347____DOLLAR__1110 =  ( n115____DOLLAR__529 ) | ( n346____DOLLAR__1109 )  ;
assign n348____DOLLAR__1111 =  ( n114____DOLLAR__525 ) | ( n347____DOLLAR__1110 )  ;
assign n349____DOLLAR__1112 =  ( n113____DOLLAR__521 ) | ( n348____DOLLAR__1111 )  ;
assign n350____DOLLAR__1113 =  ( n112____DOLLAR__517 ) | ( n349____DOLLAR__1112 )  ;
assign n351____DOLLAR__1114 =  ( n111____DOLLAR__513 ) | ( n350____DOLLAR__1113 )  ;
assign n352____DOLLAR__1115 =  ( n110____DOLLAR__509 ) | ( n351____DOLLAR__1114 )  ;
assign n353____DOLLAR__1116 =  ( n109____DOLLAR__505 ) | ( n352____DOLLAR__1115 )  ;
assign n354____DOLLAR__1117 =  ( n108____DOLLAR__501 ) | ( n353____DOLLAR__1116 )  ;
assign n355____DOLLAR__1118 =  ( n107____DOLLAR__497 ) | ( n354____DOLLAR__1117 )  ;
assign n356____DOLLAR__1119 =  ( n106____DOLLAR__493 ) | ( n355____DOLLAR__1118 )  ;
assign n357____DOLLAR__1120 =  ( n105____DOLLAR__489 ) | ( n356____DOLLAR__1119 )  ;
assign n358____DOLLAR__1121 =  ( n104____DOLLAR__485 ) | ( n357____DOLLAR__1120 )  ;
assign n359____DOLLAR__1122 =  ( n103____DOLLAR__481 ) | ( n358____DOLLAR__1121 )  ;
assign n360____DOLLAR__1123 =  ( n102____DOLLAR__477 ) | ( n359____DOLLAR__1122 )  ;
assign n361____DOLLAR__1124 =  ( n101____DOLLAR__473 ) | ( n360____DOLLAR__1123 )  ;
assign n362____DOLLAR__1125 =  ( n100____DOLLAR__469 ) | ( n361____DOLLAR__1124 )  ;
assign n363____DOLLAR__1126 =  ( n99____DOLLAR__465 ) | ( n362____DOLLAR__1125 )  ;
assign n364____DOLLAR__1127 =  ( n98____DOLLAR__461 ) | ( n363____DOLLAR__1126 )  ;
assign n365____DOLLAR__1128 =  ( n97____DOLLAR__457 ) | ( n364____DOLLAR__1127 )  ;
assign n366____DOLLAR__1129 =  ( n96____DOLLAR__453 ) | ( n365____DOLLAR__1128 )  ;
assign n367____DOLLAR__1130 =  ( n95____DOLLAR__449 ) | ( n366____DOLLAR__1129 )  ;
assign n368____DOLLAR__1131 =  ( n94____DOLLAR__445 ) | ( n367____DOLLAR__1130 )  ;
assign n369____DOLLAR__1132 =  ( n93____DOLLAR__441 ) | ( n368____DOLLAR__1131 )  ;
assign n370____DOLLAR__1133 =  ( n92____DOLLAR__437 ) | ( n369____DOLLAR__1132 )  ;
assign n371____DOLLAR__1134 =  ( n91____DOLLAR__433 ) | ( n370____DOLLAR__1133 )  ;
assign n372____DOLLAR__1135 =  ( n90____DOLLAR__429 ) | ( n371____DOLLAR__1134 )  ;
assign n373____DOLLAR__1136 =  ( n89____DOLLAR__425 ) | ( n372____DOLLAR__1135 )  ;
assign n374____DOLLAR__1137 =  ( n88____DOLLAR__421 ) | ( n373____DOLLAR__1136 )  ;
assign n375____DOLLAR__1138 =  ( n87____DOLLAR__417 ) | ( n374____DOLLAR__1137 )  ;
assign n376____DOLLAR__1139 =  ( n86____DOLLAR__413 ) | ( n375____DOLLAR__1138 )  ;
assign n377____DOLLAR__1140 =  ( n85____DOLLAR__409 ) | ( n376____DOLLAR__1139 )  ;
assign n378____DOLLAR__1141 =  ( n84____DOLLAR__405 ) | ( n377____DOLLAR__1140 )  ;
assign n379____DOLLAR__1142 =  ( n83____DOLLAR__401 ) | ( n378____DOLLAR__1141 )  ;
assign n380____DOLLAR__1143 =  ( n82____DOLLAR__397 ) | ( n379____DOLLAR__1142 )  ;
assign n381____DOLLAR__1144 =  ( n81____DOLLAR__393 ) | ( n380____DOLLAR__1143 )  ;
assign n382____DOLLAR__1145 =  ( n80____DOLLAR__389 ) | ( n381____DOLLAR__1144 )  ;
assign n383____DOLLAR__1146 =  ( n79____DOLLAR__385 ) | ( n382____DOLLAR__1145 )  ;
assign n384____DOLLAR__1147 =  ( n78____DOLLAR__381 ) | ( n383____DOLLAR__1146 )  ;
assign n385____DOLLAR__1148 =  ( n77____DOLLAR__377 ) | ( n384____DOLLAR__1147 )  ;
assign n386____DOLLAR__1149 =  ( n76____DOLLAR__373 ) | ( n385____DOLLAR__1148 )  ;
assign n387____DOLLAR__1150 =  ( n75____DOLLAR__369 ) | ( n386____DOLLAR__1149 )  ;
assign n388____DOLLAR__1151 =  ( n74____DOLLAR__365 ) | ( n387____DOLLAR__1150 )  ;
assign n389____DOLLAR__1152 =  ( n73____DOLLAR__361 ) | ( n388____DOLLAR__1151 )  ;
assign n390____DOLLAR__1153 =  ( n72____DOLLAR__357 ) | ( n389____DOLLAR__1152 )  ;
assign n391____DOLLAR__1154 =  ( n71____DOLLAR__353 ) | ( n390____DOLLAR__1153 )  ;
assign n392____DOLLAR__1155 =  ( n70____DOLLAR__349 ) | ( n391____DOLLAR__1154 )  ;
assign n393____DOLLAR__1156 =  ( n69____DOLLAR__345 ) | ( n392____DOLLAR__1155 )  ;
assign n394____DOLLAR__1157 =  ( n68____DOLLAR__341 ) | ( n393____DOLLAR__1156 )  ;
assign n395____DOLLAR__1158 =  ( n67____DOLLAR__337 ) | ( n394____DOLLAR__1157 )  ;
assign n396____DOLLAR__1159 =  ( n66____DOLLAR__333 ) | ( n395____DOLLAR__1158 )  ;
assign n397____DOLLAR__1160 =  ( n65____DOLLAR__329 ) | ( n396____DOLLAR__1159 )  ;
assign n398____DOLLAR__1161 =  ( n64____DOLLAR__325 ) | ( n397____DOLLAR__1160 )  ;
assign n399____DOLLAR__1162 =  ( n63____DOLLAR__321 ) | ( n398____DOLLAR__1161 )  ;
assign n400____DOLLAR__1163 =  ( n62____DOLLAR__317 ) | ( n399____DOLLAR__1162 )  ;
assign n401____DOLLAR__1164 =  ( n61____DOLLAR__313 ) | ( n400____DOLLAR__1163 )  ;
assign n402____DOLLAR__1165 =  ( n60____DOLLAR__309 ) | ( n401____DOLLAR__1164 )  ;
assign n403____DOLLAR__1166 =  ( n59____DOLLAR__305 ) | ( n402____DOLLAR__1165 )  ;
assign n404____DOLLAR__1167 =  ( n58____DOLLAR__301 ) | ( n403____DOLLAR__1166 )  ;
assign n405____DOLLAR__1168 =  ( n57____DOLLAR__297 ) | ( n404____DOLLAR__1167 )  ;
assign n406____DOLLAR__1169 =  ( n56____DOLLAR__293 ) | ( n405____DOLLAR__1168 )  ;
assign n407____DOLLAR__1170 =  ( n55____DOLLAR__289 ) | ( n406____DOLLAR__1169 )  ;
assign n408____DOLLAR__1171 =  ( n54____DOLLAR__285 ) | ( n407____DOLLAR__1170 )  ;
assign n409____DOLLAR__1172 =  ( n53____DOLLAR__281 ) | ( n408____DOLLAR__1171 )  ;
assign n410____DOLLAR__1173 =  ( n52____DOLLAR__277 ) | ( n409____DOLLAR__1172 )  ;
assign n411____DOLLAR__1174 =  ( n51____DOLLAR__273 ) | ( n410____DOLLAR__1173 )  ;
assign n412____DOLLAR__1175 =  ( n50____DOLLAR__269 ) | ( n411____DOLLAR__1174 )  ;
assign n413____DOLLAR__1176 =  ( n49____DOLLAR__265 ) | ( n412____DOLLAR__1175 )  ;
assign n414____DOLLAR__1177 =  ( n48____DOLLAR__261 ) | ( n413____DOLLAR__1176 )  ;
assign n415____DOLLAR__1178 =  ( n47____DOLLAR__257 ) | ( n414____DOLLAR__1177 )  ;
assign n416____DOLLAR__1179 =  ( n46____DOLLAR__253 ) | ( n415____DOLLAR__1178 )  ;
assign n417____DOLLAR__1180 =  ( n45____DOLLAR__249 ) | ( n416____DOLLAR__1179 )  ;
assign n418____DOLLAR__1181 =  ( n44____DOLLAR__245 ) | ( n417____DOLLAR__1180 )  ;
assign n419____DOLLAR__1182 =  ( n43____DOLLAR__241 ) | ( n418____DOLLAR__1181 )  ;
assign n420____DOLLAR__1183 =  ( n42____DOLLAR__237 ) | ( n419____DOLLAR__1182 )  ;
assign n421____DOLLAR__1184 =  ( n41____DOLLAR__233 ) | ( n420____DOLLAR__1183 )  ;
assign n422____DOLLAR__1185 =  ( n40____DOLLAR__229 ) | ( n421____DOLLAR__1184 )  ;
assign n423____DOLLAR__1186 =  ( n39____DOLLAR__225 ) | ( n422____DOLLAR__1185 )  ;
assign n424____DOLLAR__1187 =  ( n38____DOLLAR__221 ) | ( n423____DOLLAR__1186 )  ;
assign n425____DOLLAR__1188 =  ( n37____DOLLAR__217 ) | ( n424____DOLLAR__1187 )  ;
assign n426____DOLLAR__1189 =  ( n36____DOLLAR__213 ) | ( n425____DOLLAR__1188 )  ;
assign n427____DOLLAR__1190 =  ( n35____DOLLAR__209 ) | ( n426____DOLLAR__1189 )  ;
assign n428____DOLLAR__1191 =  ( n34____DOLLAR__205 ) | ( n427____DOLLAR__1190 )  ;
assign n429____DOLLAR__1192 =  ( n33____DOLLAR__201 ) | ( n428____DOLLAR__1191 )  ;
assign n430____DOLLAR__1193 =  ( n32____DOLLAR__197 ) | ( n429____DOLLAR__1192 )  ;
assign n431____DOLLAR__1194 =  ( n31____DOLLAR__193 ) | ( n430____DOLLAR__1193 )  ;
assign n432____DOLLAR__1195 =  ( n30____DOLLAR__189 ) | ( n431____DOLLAR__1194 )  ;
assign n433____DOLLAR__1196 =  ( n29____DOLLAR__185 ) | ( n432____DOLLAR__1195 )  ;
assign n434____DOLLAR__1197 =  ( n28____DOLLAR__181 ) | ( n433____DOLLAR__1196 )  ;
assign n435____DOLLAR__1198 =  ( n27____DOLLAR__177 ) | ( n434____DOLLAR__1197 )  ;
assign n436____DOLLAR__1199 =  ( n26____DOLLAR__173 ) | ( n435____DOLLAR__1198 )  ;
assign n437____DOLLAR__1200 =  ( n25____DOLLAR__169 ) | ( n436____DOLLAR__1199 )  ;
assign n438____DOLLAR__1201 =  ( n24____DOLLAR__165 ) | ( n437____DOLLAR__1200 )  ;
assign n439____DOLLAR__1202 =  ( n23____DOLLAR__161 ) | ( n438____DOLLAR__1201 )  ;
assign n440____DOLLAR__1203 =  ( n22____DOLLAR__157 ) | ( n439____DOLLAR__1202 )  ;
assign n441____DOLLAR__1204 =  ( n21____DOLLAR__153 ) | ( n440____DOLLAR__1203 )  ;
assign n442____DOLLAR__1205 =  ( n20____DOLLAR__149 ) | ( n441____DOLLAR__1204 )  ;
assign n443____DOLLAR__1206 =  ( n19____DOLLAR__145 ) | ( n442____DOLLAR__1205 )  ;
assign n444____DOLLAR__1207 =  ( n18____DOLLAR__141 ) | ( n443____DOLLAR__1206 )  ;
assign n445____DOLLAR__1208 =  ( n17____DOLLAR__137 ) | ( n444____DOLLAR__1207 )  ;
assign n446____DOLLAR__1209 =  ( n16____DOLLAR__133 ) | ( n445____DOLLAR__1208 )  ;
assign n447____DOLLAR__1210 =  ( n15____DOLLAR__129 ) | ( n446____DOLLAR__1209 )  ;
assign n448____DOLLAR__1211 =  ( n14____DOLLAR__125 ) | ( n447____DOLLAR__1210 )  ;
assign n449____DOLLAR__1212 =  ( n13____DOLLAR__121 ) | ( n448____DOLLAR__1211 )  ;
assign n450____DOLLAR__1213 =  ( n12____DOLLAR__117 ) | ( n449____DOLLAR__1212 )  ;
assign n451____DOLLAR__1214 =  ( n11____DOLLAR__113 ) | ( n450____DOLLAR__1213 )  ;
assign n452____DOLLAR__1215 =  ( n10____DOLLAR__109 ) | ( n451____DOLLAR__1214 )  ;
assign n453____DOLLAR__1216 =  ( n9____DOLLAR__105 ) | ( n452____DOLLAR__1215 )  ;
assign n454____DOLLAR__1217 =  ( n8____DOLLAR__101 ) | ( n453____DOLLAR__1216 )  ;
assign n455____DOLLAR__1218 =  ( n7____DOLLAR__97 ) | ( n454____DOLLAR__1217 )  ;
assign n456____DOLLAR__1219 =  ( n6____DOLLAR__93 ) | ( n455____DOLLAR__1218 )  ;
assign n457____DOLLAR__1220 =  ( n5____DOLLAR__89 ) | ( n456____DOLLAR__1219 )  ;
assign n458____DOLLAR__1221 =  ( n4____DOLLAR__85 ) | ( n457____DOLLAR__1220 )  ;
assign n459____DOLLAR__1222 =  ( n3____DOLLAR__81 ) | ( n458____DOLLAR__1221 )  ;
assign n460____DOLLAR__1223 =  ( n2____DOLLAR__77 ) | ( n459____DOLLAR__1222 )  ;
assign n461____DOLLAR__1228 =  { ( DPH ) , ( DPL ) }  ;
assign n462____DOLLAR__1230 = n461____DOLLAR__1228[7:0] ;
assign n463____DOLLAR__1232 =  ( n460____DOLLAR__1223 ) ? ( n462____DOLLAR__1230 ) : ( DPL ) ;
assign n464____DOLLAR__1237 =  ( oc8051_ROM_rdata_0 ) == ( 8'd255 )  ;
assign n465____DOLLAR__1241 =  ( oc8051_ROM_rdata_0 ) == ( 8'd254 )  ;
assign n466____DOLLAR__1245 =  ( oc8051_ROM_rdata_0 ) == ( 8'd253 )  ;
assign n467____DOLLAR__1249 =  ( oc8051_ROM_rdata_0 ) == ( 8'd252 )  ;
assign n468____DOLLAR__1253 =  ( oc8051_ROM_rdata_0 ) == ( 8'd251 )  ;
assign n469____DOLLAR__1257 =  ( oc8051_ROM_rdata_0 ) == ( 8'd250 )  ;
assign n470____DOLLAR__1261 =  ( oc8051_ROM_rdata_0 ) == ( 8'd249 )  ;
assign n471____DOLLAR__1265 =  ( oc8051_ROM_rdata_0 ) == ( 8'd248 )  ;
assign n472____DOLLAR__1269 =  ( oc8051_ROM_rdata_0 ) == ( 8'd247 )  ;
assign n473____DOLLAR__1273 =  ( oc8051_ROM_rdata_0 ) == ( 8'd246 )  ;
assign n474____DOLLAR__1277 =  ( oc8051_ROM_rdata_0 ) == ( 8'd244 )  ;
assign n475____DOLLAR__1281 =  ( oc8051_ROM_rdata_0 ) == ( 8'd243 )  ;
assign n476____DOLLAR__1285 =  ( oc8051_ROM_rdata_0 ) == ( 8'd242 )  ;
assign n477____DOLLAR__1289 =  ( oc8051_ROM_rdata_0 ) == ( 8'd241 )  ;
assign n478____DOLLAR__1293 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign n479____DOLLAR__1297 =  ( oc8051_ROM_rdata_0 ) == ( 8'd239 )  ;
assign n480____DOLLAR__1301 =  ( oc8051_ROM_rdata_0 ) == ( 8'd238 )  ;
assign n481____DOLLAR__1305 =  ( oc8051_ROM_rdata_0 ) == ( 8'd237 )  ;
assign n482____DOLLAR__1309 =  ( oc8051_ROM_rdata_0 ) == ( 8'd236 )  ;
assign n483____DOLLAR__1313 =  ( oc8051_ROM_rdata_0 ) == ( 8'd235 )  ;
assign n484____DOLLAR__1317 =  ( oc8051_ROM_rdata_0 ) == ( 8'd234 )  ;
assign n485____DOLLAR__1321 =  ( oc8051_ROM_rdata_0 ) == ( 8'd233 )  ;
assign n486____DOLLAR__1325 =  ( oc8051_ROM_rdata_0 ) == ( 8'd232 )  ;
assign n487____DOLLAR__1329 =  ( oc8051_ROM_rdata_0 ) == ( 8'd231 )  ;
assign n488____DOLLAR__1333 =  ( oc8051_ROM_rdata_0 ) == ( 8'd230 )  ;
assign n489____DOLLAR__1337 =  ( oc8051_ROM_rdata_0 ) == ( 8'd229 )  ;
assign n490____DOLLAR__1341 =  ( oc8051_ROM_rdata_0 ) == ( 8'd228 )  ;
assign n491____DOLLAR__1345 =  ( oc8051_ROM_rdata_0 ) == ( 8'd227 )  ;
assign n492____DOLLAR__1349 =  ( oc8051_ROM_rdata_0 ) == ( 8'd226 )  ;
assign n493____DOLLAR__1353 =  ( oc8051_ROM_rdata_0 ) == ( 8'd225 )  ;
assign n494____DOLLAR__1357 =  ( oc8051_ROM_rdata_0 ) == ( 8'd224 )  ;
assign n495____DOLLAR__1361 =  ( oc8051_ROM_rdata_0 ) == ( 8'd223 )  ;
assign n496____DOLLAR__1365 =  ( oc8051_ROM_rdata_0 ) == ( 8'd222 )  ;
assign n497____DOLLAR__1369 =  ( oc8051_ROM_rdata_0 ) == ( 8'd221 )  ;
assign n498____DOLLAR__1373 =  ( oc8051_ROM_rdata_0 ) == ( 8'd220 )  ;
assign n499____DOLLAR__1377 =  ( oc8051_ROM_rdata_0 ) == ( 8'd219 )  ;
assign n500____DOLLAR__1381 =  ( oc8051_ROM_rdata_0 ) == ( 8'd218 )  ;
assign n501____DOLLAR__1385 =  ( oc8051_ROM_rdata_0 ) == ( 8'd217 )  ;
assign n502____DOLLAR__1389 =  ( oc8051_ROM_rdata_0 ) == ( 8'd216 )  ;
assign n503____DOLLAR__1393 =  ( oc8051_ROM_rdata_0 ) == ( 8'd215 )  ;
assign n504____DOLLAR__1397 =  ( oc8051_ROM_rdata_0 ) == ( 8'd214 )  ;
assign n505____DOLLAR__1401 =  ( oc8051_ROM_rdata_0 ) == ( 8'd212 )  ;
assign n506____DOLLAR__1405 =  ( oc8051_ROM_rdata_0 ) == ( 8'd211 )  ;
assign n507____DOLLAR__1409 =  ( oc8051_ROM_rdata_0 ) == ( 8'd209 )  ;
assign n508____DOLLAR__1413 =  ( oc8051_ROM_rdata_0 ) == ( 8'd207 )  ;
assign n509____DOLLAR__1417 =  ( oc8051_ROM_rdata_0 ) == ( 8'd206 )  ;
assign n510____DOLLAR__1421 =  ( oc8051_ROM_rdata_0 ) == ( 8'd205 )  ;
assign n511____DOLLAR__1425 =  ( oc8051_ROM_rdata_0 ) == ( 8'd204 )  ;
assign n512____DOLLAR__1429 =  ( oc8051_ROM_rdata_0 ) == ( 8'd203 )  ;
assign n513____DOLLAR__1433 =  ( oc8051_ROM_rdata_0 ) == ( 8'd202 )  ;
assign n514____DOLLAR__1437 =  ( oc8051_ROM_rdata_0 ) == ( 8'd201 )  ;
assign n515____DOLLAR__1441 =  ( oc8051_ROM_rdata_0 ) == ( 8'd200 )  ;
assign n516____DOLLAR__1445 =  ( oc8051_ROM_rdata_0 ) == ( 8'd199 )  ;
assign n517____DOLLAR__1449 =  ( oc8051_ROM_rdata_0 ) == ( 8'd198 )  ;
assign n518____DOLLAR__1453 =  ( oc8051_ROM_rdata_0 ) == ( 8'd196 )  ;
assign n519____DOLLAR__1457 =  ( oc8051_ROM_rdata_0 ) == ( 8'd195 )  ;
assign n520____DOLLAR__1461 =  ( oc8051_ROM_rdata_0 ) == ( 8'd193 )  ;
assign n521____DOLLAR__1465 =  ( oc8051_ROM_rdata_0 ) == ( 8'd192 )  ;
assign n522____DOLLAR__1469 =  ( oc8051_ROM_rdata_0 ) == ( 8'd191 )  ;
assign n523____DOLLAR__1473 =  ( oc8051_ROM_rdata_0 ) == ( 8'd190 )  ;
assign n524____DOLLAR__1477 =  ( oc8051_ROM_rdata_0 ) == ( 8'd189 )  ;
assign n525____DOLLAR__1481 =  ( oc8051_ROM_rdata_0 ) == ( 8'd188 )  ;
assign n526____DOLLAR__1485 =  ( oc8051_ROM_rdata_0 ) == ( 8'd187 )  ;
assign n527____DOLLAR__1489 =  ( oc8051_ROM_rdata_0 ) == ( 8'd186 )  ;
assign n528____DOLLAR__1493 =  ( oc8051_ROM_rdata_0 ) == ( 8'd185 )  ;
assign n529____DOLLAR__1497 =  ( oc8051_ROM_rdata_0 ) == ( 8'd184 )  ;
assign n530____DOLLAR__1501 =  ( oc8051_ROM_rdata_0 ) == ( 8'd183 )  ;
assign n531____DOLLAR__1505 =  ( oc8051_ROM_rdata_0 ) == ( 8'd182 )  ;
assign n532____DOLLAR__1509 =  ( oc8051_ROM_rdata_0 ) == ( 8'd181 )  ;
assign n533____DOLLAR__1513 =  ( oc8051_ROM_rdata_0 ) == ( 8'd180 )  ;
assign n534____DOLLAR__1517 =  ( oc8051_ROM_rdata_0 ) == ( 8'd179 )  ;
assign n535____DOLLAR__1521 =  ( oc8051_ROM_rdata_0 ) == ( 8'd177 )  ;
assign n536____DOLLAR__1525 =  ( oc8051_ROM_rdata_0 ) == ( 8'd176 )  ;
assign n537____DOLLAR__1529 =  ( oc8051_ROM_rdata_0 ) == ( 8'd175 )  ;
assign n538____DOLLAR__1533 =  ( oc8051_ROM_rdata_0 ) == ( 8'd174 )  ;
assign n539____DOLLAR__1537 =  ( oc8051_ROM_rdata_0 ) == ( 8'd173 )  ;
assign n540____DOLLAR__1541 =  ( oc8051_ROM_rdata_0 ) == ( 8'd172 )  ;
assign n541____DOLLAR__1545 =  ( oc8051_ROM_rdata_0 ) == ( 8'd171 )  ;
assign n542____DOLLAR__1549 =  ( oc8051_ROM_rdata_0 ) == ( 8'd170 )  ;
assign n543____DOLLAR__1553 =  ( oc8051_ROM_rdata_0 ) == ( 8'd169 )  ;
assign n544____DOLLAR__1557 =  ( oc8051_ROM_rdata_0 ) == ( 8'd168 )  ;
assign n545____DOLLAR__1561 =  ( oc8051_ROM_rdata_0 ) == ( 8'd167 )  ;
assign n546____DOLLAR__1565 =  ( oc8051_ROM_rdata_0 ) == ( 8'd166 )  ;
assign n547____DOLLAR__1569 =  ( oc8051_ROM_rdata_0 ) == ( 8'd165 )  ;
assign n548____DOLLAR__1573 =  ( oc8051_ROM_rdata_0 ) == ( 8'd164 )  ;
assign n549____DOLLAR__1577 =  ( oc8051_ROM_rdata_0 ) == ( 8'd163 )  ;
assign n550____DOLLAR__1581 =  ( oc8051_ROM_rdata_0 ) == ( 8'd162 )  ;
assign n551____DOLLAR__1585 =  ( oc8051_ROM_rdata_0 ) == ( 8'd161 )  ;
assign n552____DOLLAR__1589 =  ( oc8051_ROM_rdata_0 ) == ( 8'd160 )  ;
assign n553____DOLLAR__1593 =  ( oc8051_ROM_rdata_0 ) == ( 8'd159 )  ;
assign n554____DOLLAR__1597 =  ( oc8051_ROM_rdata_0 ) == ( 8'd158 )  ;
assign n555____DOLLAR__1601 =  ( oc8051_ROM_rdata_0 ) == ( 8'd157 )  ;
assign n556____DOLLAR__1605 =  ( oc8051_ROM_rdata_0 ) == ( 8'd156 )  ;
assign n557____DOLLAR__1609 =  ( oc8051_ROM_rdata_0 ) == ( 8'd155 )  ;
assign n558____DOLLAR__1613 =  ( oc8051_ROM_rdata_0 ) == ( 8'd154 )  ;
assign n559____DOLLAR__1617 =  ( oc8051_ROM_rdata_0 ) == ( 8'd153 )  ;
assign n560____DOLLAR__1621 =  ( oc8051_ROM_rdata_0 ) == ( 8'd152 )  ;
assign n561____DOLLAR__1625 =  ( oc8051_ROM_rdata_0 ) == ( 8'd151 )  ;
assign n562____DOLLAR__1629 =  ( oc8051_ROM_rdata_0 ) == ( 8'd150 )  ;
assign n563____DOLLAR__1633 =  ( oc8051_ROM_rdata_0 ) == ( 8'd149 )  ;
assign n564____DOLLAR__1637 =  ( oc8051_ROM_rdata_0 ) == ( 8'd148 )  ;
assign n565____DOLLAR__1641 =  ( oc8051_ROM_rdata_0 ) == ( 8'd147 )  ;
assign n566____DOLLAR__1645 =  ( oc8051_ROM_rdata_0 ) == ( 8'd145 )  ;
assign n567____DOLLAR__1649 =  ( oc8051_ROM_rdata_0 ) == ( 8'd144 )  ;
assign n568____DOLLAR__1653 =  ( oc8051_ROM_rdata_0 ) == ( 8'd132 )  ;
assign n569____DOLLAR__1657 =  ( oc8051_ROM_rdata_0 ) == ( 8'd131 )  ;
assign n570____DOLLAR__1661 =  ( oc8051_ROM_rdata_0 ) == ( 8'd130 )  ;
assign n571____DOLLAR__1665 =  ( oc8051_ROM_rdata_0 ) == ( 8'd129 )  ;
assign n572____DOLLAR__1669 =  ( oc8051_ROM_rdata_0 ) == ( 8'd128 )  ;
assign n573____DOLLAR__1673 =  ( oc8051_ROM_rdata_0 ) == ( 8'd127 )  ;
assign n574____DOLLAR__1677 =  ( oc8051_ROM_rdata_0 ) == ( 8'd126 )  ;
assign n575____DOLLAR__1681 =  ( oc8051_ROM_rdata_0 ) == ( 8'd125 )  ;
assign n576____DOLLAR__1685 =  ( oc8051_ROM_rdata_0 ) == ( 8'd124 )  ;
assign n577____DOLLAR__1689 =  ( oc8051_ROM_rdata_0 ) == ( 8'd123 )  ;
assign n578____DOLLAR__1693 =  ( oc8051_ROM_rdata_0 ) == ( 8'd122 )  ;
assign n579____DOLLAR__1697 =  ( oc8051_ROM_rdata_0 ) == ( 8'd121 )  ;
assign n580____DOLLAR__1701 =  ( oc8051_ROM_rdata_0 ) == ( 8'd120 )  ;
assign n581____DOLLAR__1705 =  ( oc8051_ROM_rdata_0 ) == ( 8'd119 )  ;
assign n582____DOLLAR__1709 =  ( oc8051_ROM_rdata_0 ) == ( 8'd118 )  ;
assign n583____DOLLAR__1713 =  ( oc8051_ROM_rdata_0 ) == ( 8'd116 )  ;
assign n584____DOLLAR__1717 =  ( oc8051_ROM_rdata_0 ) == ( 8'd115 )  ;
assign n585____DOLLAR__1721 =  ( oc8051_ROM_rdata_0 ) == ( 8'd114 )  ;
assign n586____DOLLAR__1725 =  ( oc8051_ROM_rdata_0 ) == ( 8'd113 )  ;
assign n587____DOLLAR__1729 =  ( oc8051_ROM_rdata_0 ) == ( 8'd112 )  ;
assign n588____DOLLAR__1733 =  ( oc8051_ROM_rdata_0 ) == ( 8'd111 )  ;
assign n589____DOLLAR__1737 =  ( oc8051_ROM_rdata_0 ) == ( 8'd110 )  ;
assign n590____DOLLAR__1741 =  ( oc8051_ROM_rdata_0 ) == ( 8'd109 )  ;
assign n591____DOLLAR__1745 =  ( oc8051_ROM_rdata_0 ) == ( 8'd108 )  ;
assign n592____DOLLAR__1749 =  ( oc8051_ROM_rdata_0 ) == ( 8'd107 )  ;
assign n593____DOLLAR__1753 =  ( oc8051_ROM_rdata_0 ) == ( 8'd106 )  ;
assign n594____DOLLAR__1757 =  ( oc8051_ROM_rdata_0 ) == ( 8'd105 )  ;
assign n595____DOLLAR__1761 =  ( oc8051_ROM_rdata_0 ) == ( 8'd104 )  ;
assign n596____DOLLAR__1765 =  ( oc8051_ROM_rdata_0 ) == ( 8'd103 )  ;
assign n597____DOLLAR__1769 =  ( oc8051_ROM_rdata_0 ) == ( 8'd102 )  ;
assign n598____DOLLAR__1773 =  ( oc8051_ROM_rdata_0 ) == ( 8'd101 )  ;
assign n599____DOLLAR__1777 =  ( oc8051_ROM_rdata_0 ) == ( 8'd100 )  ;
assign n600____DOLLAR__1781 =  ( oc8051_ROM_rdata_0 ) == ( 8'd97 )  ;
assign n601____DOLLAR__1785 =  ( oc8051_ROM_rdata_0 ) == ( 8'd96 )  ;
assign n602____DOLLAR__1789 =  ( oc8051_ROM_rdata_0 ) == ( 8'd95 )  ;
assign n603____DOLLAR__1793 =  ( oc8051_ROM_rdata_0 ) == ( 8'd94 )  ;
assign n604____DOLLAR__1797 =  ( oc8051_ROM_rdata_0 ) == ( 8'd93 )  ;
assign n605____DOLLAR__1801 =  ( oc8051_ROM_rdata_0 ) == ( 8'd92 )  ;
assign n606____DOLLAR__1805 =  ( oc8051_ROM_rdata_0 ) == ( 8'd91 )  ;
assign n607____DOLLAR__1809 =  ( oc8051_ROM_rdata_0 ) == ( 8'd90 )  ;
assign n608____DOLLAR__1813 =  ( oc8051_ROM_rdata_0 ) == ( 8'd89 )  ;
assign n609____DOLLAR__1817 =  ( oc8051_ROM_rdata_0 ) == ( 8'd88 )  ;
assign n610____DOLLAR__1821 =  ( oc8051_ROM_rdata_0 ) == ( 8'd87 )  ;
assign n611____DOLLAR__1825 =  ( oc8051_ROM_rdata_0 ) == ( 8'd86 )  ;
assign n612____DOLLAR__1829 =  ( oc8051_ROM_rdata_0 ) == ( 8'd85 )  ;
assign n613____DOLLAR__1833 =  ( oc8051_ROM_rdata_0 ) == ( 8'd84 )  ;
assign n614____DOLLAR__1837 =  ( oc8051_ROM_rdata_0 ) == ( 8'd81 )  ;
assign n615____DOLLAR__1841 =  ( oc8051_ROM_rdata_0 ) == ( 8'd80 )  ;
assign n616____DOLLAR__1845 =  ( oc8051_ROM_rdata_0 ) == ( 8'd79 )  ;
assign n617____DOLLAR__1849 =  ( oc8051_ROM_rdata_0 ) == ( 8'd78 )  ;
assign n618____DOLLAR__1853 =  ( oc8051_ROM_rdata_0 ) == ( 8'd77 )  ;
assign n619____DOLLAR__1857 =  ( oc8051_ROM_rdata_0 ) == ( 8'd76 )  ;
assign n620____DOLLAR__1861 =  ( oc8051_ROM_rdata_0 ) == ( 8'd75 )  ;
assign n621____DOLLAR__1865 =  ( oc8051_ROM_rdata_0 ) == ( 8'd74 )  ;
assign n622____DOLLAR__1869 =  ( oc8051_ROM_rdata_0 ) == ( 8'd73 )  ;
assign n623____DOLLAR__1873 =  ( oc8051_ROM_rdata_0 ) == ( 8'd72 )  ;
assign n624____DOLLAR__1877 =  ( oc8051_ROM_rdata_0 ) == ( 8'd71 )  ;
assign n625____DOLLAR__1881 =  ( oc8051_ROM_rdata_0 ) == ( 8'd70 )  ;
assign n626____DOLLAR__1885 =  ( oc8051_ROM_rdata_0 ) == ( 8'd69 )  ;
assign n627____DOLLAR__1889 =  ( oc8051_ROM_rdata_0 ) == ( 8'd68 )  ;
assign n628____DOLLAR__1893 =  ( oc8051_ROM_rdata_0 ) == ( 8'd65 )  ;
assign n629____DOLLAR__1897 =  ( oc8051_ROM_rdata_0 ) == ( 8'd64 )  ;
assign n630____DOLLAR__1901 =  ( oc8051_ROM_rdata_0 ) == ( 8'd63 )  ;
assign n631____DOLLAR__1905 =  ( oc8051_ROM_rdata_0 ) == ( 8'd62 )  ;
assign n632____DOLLAR__1909 =  ( oc8051_ROM_rdata_0 ) == ( 8'd61 )  ;
assign n633____DOLLAR__1913 =  ( oc8051_ROM_rdata_0 ) == ( 8'd60 )  ;
assign n634____DOLLAR__1917 =  ( oc8051_ROM_rdata_0 ) == ( 8'd59 )  ;
assign n635____DOLLAR__1921 =  ( oc8051_ROM_rdata_0 ) == ( 8'd58 )  ;
assign n636____DOLLAR__1925 =  ( oc8051_ROM_rdata_0 ) == ( 8'd57 )  ;
assign n637____DOLLAR__1929 =  ( oc8051_ROM_rdata_0 ) == ( 8'd56 )  ;
assign n638____DOLLAR__1933 =  ( oc8051_ROM_rdata_0 ) == ( 8'd55 )  ;
assign n639____DOLLAR__1937 =  ( oc8051_ROM_rdata_0 ) == ( 8'd54 )  ;
assign n640____DOLLAR__1941 =  ( oc8051_ROM_rdata_0 ) == ( 8'd53 )  ;
assign n641____DOLLAR__1945 =  ( oc8051_ROM_rdata_0 ) == ( 8'd52 )  ;
assign n642____DOLLAR__1949 =  ( oc8051_ROM_rdata_0 ) == ( 8'd51 )  ;
assign n643____DOLLAR__1953 =  ( oc8051_ROM_rdata_0 ) == ( 8'd50 )  ;
assign n644____DOLLAR__1957 =  ( oc8051_ROM_rdata_0 ) == ( 8'd49 )  ;
assign n645____DOLLAR__1961 =  ( oc8051_ROM_rdata_0 ) == ( 8'd48 )  ;
assign n646____DOLLAR__1965 =  ( oc8051_ROM_rdata_0 ) == ( 8'd47 )  ;
assign n647____DOLLAR__1969 =  ( oc8051_ROM_rdata_0 ) == ( 8'd46 )  ;
assign n648____DOLLAR__1973 =  ( oc8051_ROM_rdata_0 ) == ( 8'd45 )  ;
assign n649____DOLLAR__1977 =  ( oc8051_ROM_rdata_0 ) == ( 8'd44 )  ;
assign n650____DOLLAR__1981 =  ( oc8051_ROM_rdata_0 ) == ( 8'd43 )  ;
assign n651____DOLLAR__1985 =  ( oc8051_ROM_rdata_0 ) == ( 8'd42 )  ;
assign n652____DOLLAR__1989 =  ( oc8051_ROM_rdata_0 ) == ( 8'd41 )  ;
assign n653____DOLLAR__1993 =  ( oc8051_ROM_rdata_0 ) == ( 8'd40 )  ;
assign n654____DOLLAR__1997 =  ( oc8051_ROM_rdata_0 ) == ( 8'd39 )  ;
assign n655____DOLLAR__2001 =  ( oc8051_ROM_rdata_0 ) == ( 8'd38 )  ;
assign n656____DOLLAR__2005 =  ( oc8051_ROM_rdata_0 ) == ( 8'd37 )  ;
assign n657____DOLLAR__2009 =  ( oc8051_ROM_rdata_0 ) == ( 8'd36 )  ;
assign n658____DOLLAR__2013 =  ( oc8051_ROM_rdata_0 ) == ( 8'd35 )  ;
assign n659____DOLLAR__2017 =  ( oc8051_ROM_rdata_0 ) == ( 8'd34 )  ;
assign n660____DOLLAR__2021 =  ( oc8051_ROM_rdata_0 ) == ( 8'd33 )  ;
assign n661____DOLLAR__2025 =  ( oc8051_ROM_rdata_0 ) == ( 8'd32 )  ;
assign n662____DOLLAR__2029 =  ( oc8051_ROM_rdata_0 ) == ( 8'd31 )  ;
assign n663____DOLLAR__2033 =  ( oc8051_ROM_rdata_0 ) == ( 8'd30 )  ;
assign n664____DOLLAR__2037 =  ( oc8051_ROM_rdata_0 ) == ( 8'd29 )  ;
assign n665____DOLLAR__2041 =  ( oc8051_ROM_rdata_0 ) == ( 8'd28 )  ;
assign n666____DOLLAR__2045 =  ( oc8051_ROM_rdata_0 ) == ( 8'd27 )  ;
assign n667____DOLLAR__2049 =  ( oc8051_ROM_rdata_0 ) == ( 8'd26 )  ;
assign n668____DOLLAR__2053 =  ( oc8051_ROM_rdata_0 ) == ( 8'd25 )  ;
assign n669____DOLLAR__2057 =  ( oc8051_ROM_rdata_0 ) == ( 8'd24 )  ;
assign n670____DOLLAR__2061 =  ( oc8051_ROM_rdata_0 ) == ( 8'd23 )  ;
assign n671____DOLLAR__2065 =  ( oc8051_ROM_rdata_0 ) == ( 8'd22 )  ;
assign n672____DOLLAR__2069 =  ( oc8051_ROM_rdata_0 ) == ( 8'd20 )  ;
assign n673____DOLLAR__2073 =  ( oc8051_ROM_rdata_0 ) == ( 8'd19 )  ;
assign n674____DOLLAR__2077 =  ( oc8051_ROM_rdata_0 ) == ( 8'd18 )  ;
assign n675____DOLLAR__2081 =  ( oc8051_ROM_rdata_0 ) == ( 8'd17 )  ;
assign n676____DOLLAR__2085 =  ( oc8051_ROM_rdata_0 ) == ( 8'd15 )  ;
assign n677____DOLLAR__2089 =  ( oc8051_ROM_rdata_0 ) == ( 8'd14 )  ;
assign n678____DOLLAR__2093 =  ( oc8051_ROM_rdata_0 ) == ( 8'd13 )  ;
assign n679____DOLLAR__2097 =  ( oc8051_ROM_rdata_0 ) == ( 8'd12 )  ;
assign n680____DOLLAR__2101 =  ( oc8051_ROM_rdata_0 ) == ( 8'd11 )  ;
assign n681____DOLLAR__2105 =  ( oc8051_ROM_rdata_0 ) == ( 8'd10 )  ;
assign n682____DOLLAR__2109 =  ( oc8051_ROM_rdata_0 ) == ( 8'd9 )  ;
assign n683____DOLLAR__2113 =  ( oc8051_ROM_rdata_0 ) == ( 8'd8 )  ;
assign n684____DOLLAR__2117 =  ( oc8051_ROM_rdata_0 ) == ( 8'd7 )  ;
assign n685____DOLLAR__2121 =  ( oc8051_ROM_rdata_0 ) == ( 8'd6 )  ;
assign n686____DOLLAR__2125 =  ( oc8051_ROM_rdata_0 ) == ( 8'd4 )  ;
assign n687____DOLLAR__2129 =  ( oc8051_ROM_rdata_0 ) == ( 8'd3 )  ;
assign n688____DOLLAR__2133 =  ( oc8051_ROM_rdata_0 ) == ( 8'd2 )  ;
assign n689____DOLLAR__2137 =  ( oc8051_ROM_rdata_0 ) == ( 8'd1 )  ;
assign n690____DOLLAR__2141 =  ( oc8051_ROM_rdata_0 ) == ( 8'd0 )  ;
assign n691____DOLLAR__2143 =  ( n689____DOLLAR__2137 ) | ( n690____DOLLAR__2141 )  ;
assign n692____DOLLAR__2144 =  ( n688____DOLLAR__2133 ) | ( n691____DOLLAR__2143 )  ;
assign n693____DOLLAR__2145 =  ( n687____DOLLAR__2129 ) | ( n692____DOLLAR__2144 )  ;
assign n694____DOLLAR__2146 =  ( n686____DOLLAR__2125 ) | ( n693____DOLLAR__2145 )  ;
assign n695____DOLLAR__2147 =  ( n685____DOLLAR__2121 ) | ( n694____DOLLAR__2146 )  ;
assign n696____DOLLAR__2148 =  ( n684____DOLLAR__2117 ) | ( n695____DOLLAR__2147 )  ;
assign n697____DOLLAR__2149 =  ( n683____DOLLAR__2113 ) | ( n696____DOLLAR__2148 )  ;
assign n698____DOLLAR__2150 =  ( n682____DOLLAR__2109 ) | ( n697____DOLLAR__2149 )  ;
assign n699____DOLLAR__2151 =  ( n681____DOLLAR__2105 ) | ( n698____DOLLAR__2150 )  ;
assign n700____DOLLAR__2152 =  ( n680____DOLLAR__2101 ) | ( n699____DOLLAR__2151 )  ;
assign n701____DOLLAR__2153 =  ( n679____DOLLAR__2097 ) | ( n700____DOLLAR__2152 )  ;
assign n702____DOLLAR__2154 =  ( n678____DOLLAR__2093 ) | ( n701____DOLLAR__2153 )  ;
assign n703____DOLLAR__2155 =  ( n677____DOLLAR__2089 ) | ( n702____DOLLAR__2154 )  ;
assign n704____DOLLAR__2156 =  ( n676____DOLLAR__2085 ) | ( n703____DOLLAR__2155 )  ;
assign n705____DOLLAR__2157 =  ( n675____DOLLAR__2081 ) | ( n704____DOLLAR__2156 )  ;
assign n706____DOLLAR__2158 =  ( n674____DOLLAR__2077 ) | ( n705____DOLLAR__2157 )  ;
assign n707____DOLLAR__2159 =  ( n673____DOLLAR__2073 ) | ( n706____DOLLAR__2158 )  ;
assign n708____DOLLAR__2160 =  ( n672____DOLLAR__2069 ) | ( n707____DOLLAR__2159 )  ;
assign n709____DOLLAR__2161 =  ( n671____DOLLAR__2065 ) | ( n708____DOLLAR__2160 )  ;
assign n710____DOLLAR__2162 =  ( n670____DOLLAR__2061 ) | ( n709____DOLLAR__2161 )  ;
assign n711____DOLLAR__2163 =  ( n669____DOLLAR__2057 ) | ( n710____DOLLAR__2162 )  ;
assign n712____DOLLAR__2164 =  ( n668____DOLLAR__2053 ) | ( n711____DOLLAR__2163 )  ;
assign n713____DOLLAR__2165 =  ( n667____DOLLAR__2049 ) | ( n712____DOLLAR__2164 )  ;
assign n714____DOLLAR__2166 =  ( n666____DOLLAR__2045 ) | ( n713____DOLLAR__2165 )  ;
assign n715____DOLLAR__2167 =  ( n665____DOLLAR__2041 ) | ( n714____DOLLAR__2166 )  ;
assign n716____DOLLAR__2168 =  ( n664____DOLLAR__2037 ) | ( n715____DOLLAR__2167 )  ;
assign n717____DOLLAR__2169 =  ( n663____DOLLAR__2033 ) | ( n716____DOLLAR__2168 )  ;
assign n718____DOLLAR__2170 =  ( n662____DOLLAR__2029 ) | ( n717____DOLLAR__2169 )  ;
assign n719____DOLLAR__2171 =  ( n661____DOLLAR__2025 ) | ( n718____DOLLAR__2170 )  ;
assign n720____DOLLAR__2172 =  ( n660____DOLLAR__2021 ) | ( n719____DOLLAR__2171 )  ;
assign n721____DOLLAR__2173 =  ( n659____DOLLAR__2017 ) | ( n720____DOLLAR__2172 )  ;
assign n722____DOLLAR__2174 =  ( n658____DOLLAR__2013 ) | ( n721____DOLLAR__2173 )  ;
assign n723____DOLLAR__2175 =  ( n657____DOLLAR__2009 ) | ( n722____DOLLAR__2174 )  ;
assign n724____DOLLAR__2176 =  ( n656____DOLLAR__2005 ) | ( n723____DOLLAR__2175 )  ;
assign n725____DOLLAR__2177 =  ( n655____DOLLAR__2001 ) | ( n724____DOLLAR__2176 )  ;
assign n726____DOLLAR__2178 =  ( n654____DOLLAR__1997 ) | ( n725____DOLLAR__2177 )  ;
assign n727____DOLLAR__2179 =  ( n653____DOLLAR__1993 ) | ( n726____DOLLAR__2178 )  ;
assign n728____DOLLAR__2180 =  ( n652____DOLLAR__1989 ) | ( n727____DOLLAR__2179 )  ;
assign n729____DOLLAR__2181 =  ( n651____DOLLAR__1985 ) | ( n728____DOLLAR__2180 )  ;
assign n730____DOLLAR__2182 =  ( n650____DOLLAR__1981 ) | ( n729____DOLLAR__2181 )  ;
assign n731____DOLLAR__2183 =  ( n649____DOLLAR__1977 ) | ( n730____DOLLAR__2182 )  ;
assign n732____DOLLAR__2184 =  ( n648____DOLLAR__1973 ) | ( n731____DOLLAR__2183 )  ;
assign n733____DOLLAR__2185 =  ( n647____DOLLAR__1969 ) | ( n732____DOLLAR__2184 )  ;
assign n734____DOLLAR__2186 =  ( n646____DOLLAR__1965 ) | ( n733____DOLLAR__2185 )  ;
assign n735____DOLLAR__2187 =  ( n645____DOLLAR__1961 ) | ( n734____DOLLAR__2186 )  ;
assign n736____DOLLAR__2188 =  ( n644____DOLLAR__1957 ) | ( n735____DOLLAR__2187 )  ;
assign n737____DOLLAR__2189 =  ( n643____DOLLAR__1953 ) | ( n736____DOLLAR__2188 )  ;
assign n738____DOLLAR__2190 =  ( n642____DOLLAR__1949 ) | ( n737____DOLLAR__2189 )  ;
assign n739____DOLLAR__2191 =  ( n641____DOLLAR__1945 ) | ( n738____DOLLAR__2190 )  ;
assign n740____DOLLAR__2192 =  ( n640____DOLLAR__1941 ) | ( n739____DOLLAR__2191 )  ;
assign n741____DOLLAR__2193 =  ( n639____DOLLAR__1937 ) | ( n740____DOLLAR__2192 )  ;
assign n742____DOLLAR__2194 =  ( n638____DOLLAR__1933 ) | ( n741____DOLLAR__2193 )  ;
assign n743____DOLLAR__2195 =  ( n637____DOLLAR__1929 ) | ( n742____DOLLAR__2194 )  ;
assign n744____DOLLAR__2196 =  ( n636____DOLLAR__1925 ) | ( n743____DOLLAR__2195 )  ;
assign n745____DOLLAR__2197 =  ( n635____DOLLAR__1921 ) | ( n744____DOLLAR__2196 )  ;
assign n746____DOLLAR__2198 =  ( n634____DOLLAR__1917 ) | ( n745____DOLLAR__2197 )  ;
assign n747____DOLLAR__2199 =  ( n633____DOLLAR__1913 ) | ( n746____DOLLAR__2198 )  ;
assign n748____DOLLAR__2200 =  ( n632____DOLLAR__1909 ) | ( n747____DOLLAR__2199 )  ;
assign n749____DOLLAR__2201 =  ( n631____DOLLAR__1905 ) | ( n748____DOLLAR__2200 )  ;
assign n750____DOLLAR__2202 =  ( n630____DOLLAR__1901 ) | ( n749____DOLLAR__2201 )  ;
assign n751____DOLLAR__2203 =  ( n629____DOLLAR__1897 ) | ( n750____DOLLAR__2202 )  ;
assign n752____DOLLAR__2204 =  ( n628____DOLLAR__1893 ) | ( n751____DOLLAR__2203 )  ;
assign n753____DOLLAR__2205 =  ( n627____DOLLAR__1889 ) | ( n752____DOLLAR__2204 )  ;
assign n754____DOLLAR__2206 =  ( n626____DOLLAR__1885 ) | ( n753____DOLLAR__2205 )  ;
assign n755____DOLLAR__2207 =  ( n625____DOLLAR__1881 ) | ( n754____DOLLAR__2206 )  ;
assign n756____DOLLAR__2208 =  ( n624____DOLLAR__1877 ) | ( n755____DOLLAR__2207 )  ;
assign n757____DOLLAR__2209 =  ( n623____DOLLAR__1873 ) | ( n756____DOLLAR__2208 )  ;
assign n758____DOLLAR__2210 =  ( n622____DOLLAR__1869 ) | ( n757____DOLLAR__2209 )  ;
assign n759____DOLLAR__2211 =  ( n621____DOLLAR__1865 ) | ( n758____DOLLAR__2210 )  ;
assign n760____DOLLAR__2212 =  ( n620____DOLLAR__1861 ) | ( n759____DOLLAR__2211 )  ;
assign n761____DOLLAR__2213 =  ( n619____DOLLAR__1857 ) | ( n760____DOLLAR__2212 )  ;
assign n762____DOLLAR__2214 =  ( n618____DOLLAR__1853 ) | ( n761____DOLLAR__2213 )  ;
assign n763____DOLLAR__2215 =  ( n617____DOLLAR__1849 ) | ( n762____DOLLAR__2214 )  ;
assign n764____DOLLAR__2216 =  ( n616____DOLLAR__1845 ) | ( n763____DOLLAR__2215 )  ;
assign n765____DOLLAR__2217 =  ( n615____DOLLAR__1841 ) | ( n764____DOLLAR__2216 )  ;
assign n766____DOLLAR__2218 =  ( n614____DOLLAR__1837 ) | ( n765____DOLLAR__2217 )  ;
assign n767____DOLLAR__2219 =  ( n613____DOLLAR__1833 ) | ( n766____DOLLAR__2218 )  ;
assign n768____DOLLAR__2220 =  ( n612____DOLLAR__1829 ) | ( n767____DOLLAR__2219 )  ;
assign n769____DOLLAR__2221 =  ( n611____DOLLAR__1825 ) | ( n768____DOLLAR__2220 )  ;
assign n770____DOLLAR__2222 =  ( n610____DOLLAR__1821 ) | ( n769____DOLLAR__2221 )  ;
assign n771____DOLLAR__2223 =  ( n609____DOLLAR__1817 ) | ( n770____DOLLAR__2222 )  ;
assign n772____DOLLAR__2224 =  ( n608____DOLLAR__1813 ) | ( n771____DOLLAR__2223 )  ;
assign n773____DOLLAR__2225 =  ( n607____DOLLAR__1809 ) | ( n772____DOLLAR__2224 )  ;
assign n774____DOLLAR__2226 =  ( n606____DOLLAR__1805 ) | ( n773____DOLLAR__2225 )  ;
assign n775____DOLLAR__2227 =  ( n605____DOLLAR__1801 ) | ( n774____DOLLAR__2226 )  ;
assign n776____DOLLAR__2228 =  ( n604____DOLLAR__1797 ) | ( n775____DOLLAR__2227 )  ;
assign n777____DOLLAR__2229 =  ( n603____DOLLAR__1793 ) | ( n776____DOLLAR__2228 )  ;
assign n778____DOLLAR__2230 =  ( n602____DOLLAR__1789 ) | ( n777____DOLLAR__2229 )  ;
assign n779____DOLLAR__2231 =  ( n601____DOLLAR__1785 ) | ( n778____DOLLAR__2230 )  ;
assign n780____DOLLAR__2232 =  ( n600____DOLLAR__1781 ) | ( n779____DOLLAR__2231 )  ;
assign n781____DOLLAR__2233 =  ( n599____DOLLAR__1777 ) | ( n780____DOLLAR__2232 )  ;
assign n782____DOLLAR__2234 =  ( n598____DOLLAR__1773 ) | ( n781____DOLLAR__2233 )  ;
assign n783____DOLLAR__2235 =  ( n597____DOLLAR__1769 ) | ( n782____DOLLAR__2234 )  ;
assign n784____DOLLAR__2236 =  ( n596____DOLLAR__1765 ) | ( n783____DOLLAR__2235 )  ;
assign n785____DOLLAR__2237 =  ( n595____DOLLAR__1761 ) | ( n784____DOLLAR__2236 )  ;
assign n786____DOLLAR__2238 =  ( n594____DOLLAR__1757 ) | ( n785____DOLLAR__2237 )  ;
assign n787____DOLLAR__2239 =  ( n593____DOLLAR__1753 ) | ( n786____DOLLAR__2238 )  ;
assign n788____DOLLAR__2240 =  ( n592____DOLLAR__1749 ) | ( n787____DOLLAR__2239 )  ;
assign n789____DOLLAR__2241 =  ( n591____DOLLAR__1745 ) | ( n788____DOLLAR__2240 )  ;
assign n790____DOLLAR__2242 =  ( n590____DOLLAR__1741 ) | ( n789____DOLLAR__2241 )  ;
assign n791____DOLLAR__2243 =  ( n589____DOLLAR__1737 ) | ( n790____DOLLAR__2242 )  ;
assign n792____DOLLAR__2244 =  ( n588____DOLLAR__1733 ) | ( n791____DOLLAR__2243 )  ;
assign n793____DOLLAR__2245 =  ( n587____DOLLAR__1729 ) | ( n792____DOLLAR__2244 )  ;
assign n794____DOLLAR__2246 =  ( n586____DOLLAR__1725 ) | ( n793____DOLLAR__2245 )  ;
assign n795____DOLLAR__2247 =  ( n585____DOLLAR__1721 ) | ( n794____DOLLAR__2246 )  ;
assign n796____DOLLAR__2248 =  ( n584____DOLLAR__1717 ) | ( n795____DOLLAR__2247 )  ;
assign n797____DOLLAR__2249 =  ( n583____DOLLAR__1713 ) | ( n796____DOLLAR__2248 )  ;
assign n798____DOLLAR__2250 =  ( n582____DOLLAR__1709 ) | ( n797____DOLLAR__2249 )  ;
assign n799____DOLLAR__2251 =  ( n581____DOLLAR__1705 ) | ( n798____DOLLAR__2250 )  ;
assign n800____DOLLAR__2252 =  ( n580____DOLLAR__1701 ) | ( n799____DOLLAR__2251 )  ;
assign n801____DOLLAR__2253 =  ( n579____DOLLAR__1697 ) | ( n800____DOLLAR__2252 )  ;
assign n802____DOLLAR__2254 =  ( n578____DOLLAR__1693 ) | ( n801____DOLLAR__2253 )  ;
assign n803____DOLLAR__2255 =  ( n577____DOLLAR__1689 ) | ( n802____DOLLAR__2254 )  ;
assign n804____DOLLAR__2256 =  ( n576____DOLLAR__1685 ) | ( n803____DOLLAR__2255 )  ;
assign n805____DOLLAR__2257 =  ( n575____DOLLAR__1681 ) | ( n804____DOLLAR__2256 )  ;
assign n806____DOLLAR__2258 =  ( n574____DOLLAR__1677 ) | ( n805____DOLLAR__2257 )  ;
assign n807____DOLLAR__2259 =  ( n573____DOLLAR__1673 ) | ( n806____DOLLAR__2258 )  ;
assign n808____DOLLAR__2260 =  ( n572____DOLLAR__1669 ) | ( n807____DOLLAR__2259 )  ;
assign n809____DOLLAR__2261 =  ( n571____DOLLAR__1665 ) | ( n808____DOLLAR__2260 )  ;
assign n810____DOLLAR__2262 =  ( n570____DOLLAR__1661 ) | ( n809____DOLLAR__2261 )  ;
assign n811____DOLLAR__2263 =  ( n569____DOLLAR__1657 ) | ( n810____DOLLAR__2262 )  ;
assign n812____DOLLAR__2264 =  ( n568____DOLLAR__1653 ) | ( n811____DOLLAR__2263 )  ;
assign n813____DOLLAR__2265 =  ( n567____DOLLAR__1649 ) | ( n812____DOLLAR__2264 )  ;
assign n814____DOLLAR__2266 =  ( n566____DOLLAR__1645 ) | ( n813____DOLLAR__2265 )  ;
assign n815____DOLLAR__2267 =  ( n565____DOLLAR__1641 ) | ( n814____DOLLAR__2266 )  ;
assign n816____DOLLAR__2268 =  ( n564____DOLLAR__1637 ) | ( n815____DOLLAR__2267 )  ;
assign n817____DOLLAR__2269 =  ( n563____DOLLAR__1633 ) | ( n816____DOLLAR__2268 )  ;
assign n818____DOLLAR__2270 =  ( n562____DOLLAR__1629 ) | ( n817____DOLLAR__2269 )  ;
assign n819____DOLLAR__2271 =  ( n561____DOLLAR__1625 ) | ( n818____DOLLAR__2270 )  ;
assign n820____DOLLAR__2272 =  ( n560____DOLLAR__1621 ) | ( n819____DOLLAR__2271 )  ;
assign n821____DOLLAR__2273 =  ( n559____DOLLAR__1617 ) | ( n820____DOLLAR__2272 )  ;
assign n822____DOLLAR__2274 =  ( n558____DOLLAR__1613 ) | ( n821____DOLLAR__2273 )  ;
assign n823____DOLLAR__2275 =  ( n557____DOLLAR__1609 ) | ( n822____DOLLAR__2274 )  ;
assign n824____DOLLAR__2276 =  ( n556____DOLLAR__1605 ) | ( n823____DOLLAR__2275 )  ;
assign n825____DOLLAR__2277 =  ( n555____DOLLAR__1601 ) | ( n824____DOLLAR__2276 )  ;
assign n826____DOLLAR__2278 =  ( n554____DOLLAR__1597 ) | ( n825____DOLLAR__2277 )  ;
assign n827____DOLLAR__2279 =  ( n553____DOLLAR__1593 ) | ( n826____DOLLAR__2278 )  ;
assign n828____DOLLAR__2280 =  ( n552____DOLLAR__1589 ) | ( n827____DOLLAR__2279 )  ;
assign n829____DOLLAR__2281 =  ( n551____DOLLAR__1585 ) | ( n828____DOLLAR__2280 )  ;
assign n830____DOLLAR__2282 =  ( n550____DOLLAR__1581 ) | ( n829____DOLLAR__2281 )  ;
assign n831____DOLLAR__2283 =  ( n549____DOLLAR__1577 ) | ( n830____DOLLAR__2282 )  ;
assign n832____DOLLAR__2284 =  ( n548____DOLLAR__1573 ) | ( n831____DOLLAR__2283 )  ;
assign n833____DOLLAR__2285 =  ( n547____DOLLAR__1569 ) | ( n832____DOLLAR__2284 )  ;
assign n834____DOLLAR__2286 =  ( n546____DOLLAR__1565 ) | ( n833____DOLLAR__2285 )  ;
assign n835____DOLLAR__2287 =  ( n545____DOLLAR__1561 ) | ( n834____DOLLAR__2286 )  ;
assign n836____DOLLAR__2288 =  ( n544____DOLLAR__1557 ) | ( n835____DOLLAR__2287 )  ;
assign n837____DOLLAR__2289 =  ( n543____DOLLAR__1553 ) | ( n836____DOLLAR__2288 )  ;
assign n838____DOLLAR__2290 =  ( n542____DOLLAR__1549 ) | ( n837____DOLLAR__2289 )  ;
assign n839____DOLLAR__2291 =  ( n541____DOLLAR__1545 ) | ( n838____DOLLAR__2290 )  ;
assign n840____DOLLAR__2292 =  ( n540____DOLLAR__1541 ) | ( n839____DOLLAR__2291 )  ;
assign n841____DOLLAR__2293 =  ( n539____DOLLAR__1537 ) | ( n840____DOLLAR__2292 )  ;
assign n842____DOLLAR__2294 =  ( n538____DOLLAR__1533 ) | ( n841____DOLLAR__2293 )  ;
assign n843____DOLLAR__2295 =  ( n537____DOLLAR__1529 ) | ( n842____DOLLAR__2294 )  ;
assign n844____DOLLAR__2296 =  ( n536____DOLLAR__1525 ) | ( n843____DOLLAR__2295 )  ;
assign n845____DOLLAR__2297 =  ( n535____DOLLAR__1521 ) | ( n844____DOLLAR__2296 )  ;
assign n846____DOLLAR__2298 =  ( n534____DOLLAR__1517 ) | ( n845____DOLLAR__2297 )  ;
assign n847____DOLLAR__2299 =  ( n533____DOLLAR__1513 ) | ( n846____DOLLAR__2298 )  ;
assign n848____DOLLAR__2300 =  ( n532____DOLLAR__1509 ) | ( n847____DOLLAR__2299 )  ;
assign n849____DOLLAR__2301 =  ( n531____DOLLAR__1505 ) | ( n848____DOLLAR__2300 )  ;
assign n850____DOLLAR__2302 =  ( n530____DOLLAR__1501 ) | ( n849____DOLLAR__2301 )  ;
assign n851____DOLLAR__2303 =  ( n529____DOLLAR__1497 ) | ( n850____DOLLAR__2302 )  ;
assign n852____DOLLAR__2304 =  ( n528____DOLLAR__1493 ) | ( n851____DOLLAR__2303 )  ;
assign n853____DOLLAR__2305 =  ( n527____DOLLAR__1489 ) | ( n852____DOLLAR__2304 )  ;
assign n854____DOLLAR__2306 =  ( n526____DOLLAR__1485 ) | ( n853____DOLLAR__2305 )  ;
assign n855____DOLLAR__2307 =  ( n525____DOLLAR__1481 ) | ( n854____DOLLAR__2306 )  ;
assign n856____DOLLAR__2308 =  ( n524____DOLLAR__1477 ) | ( n855____DOLLAR__2307 )  ;
assign n857____DOLLAR__2309 =  ( n523____DOLLAR__1473 ) | ( n856____DOLLAR__2308 )  ;
assign n858____DOLLAR__2310 =  ( n522____DOLLAR__1469 ) | ( n857____DOLLAR__2309 )  ;
assign n859____DOLLAR__2311 =  ( n521____DOLLAR__1465 ) | ( n858____DOLLAR__2310 )  ;
assign n860____DOLLAR__2312 =  ( n520____DOLLAR__1461 ) | ( n859____DOLLAR__2311 )  ;
assign n861____DOLLAR__2313 =  ( n519____DOLLAR__1457 ) | ( n860____DOLLAR__2312 )  ;
assign n862____DOLLAR__2314 =  ( n518____DOLLAR__1453 ) | ( n861____DOLLAR__2313 )  ;
assign n863____DOLLAR__2315 =  ( n517____DOLLAR__1449 ) | ( n862____DOLLAR__2314 )  ;
assign n864____DOLLAR__2316 =  ( n516____DOLLAR__1445 ) | ( n863____DOLLAR__2315 )  ;
assign n865____DOLLAR__2317 =  ( n515____DOLLAR__1441 ) | ( n864____DOLLAR__2316 )  ;
assign n866____DOLLAR__2318 =  ( n514____DOLLAR__1437 ) | ( n865____DOLLAR__2317 )  ;
assign n867____DOLLAR__2319 =  ( n513____DOLLAR__1433 ) | ( n866____DOLLAR__2318 )  ;
assign n868____DOLLAR__2320 =  ( n512____DOLLAR__1429 ) | ( n867____DOLLAR__2319 )  ;
assign n869____DOLLAR__2321 =  ( n511____DOLLAR__1425 ) | ( n868____DOLLAR__2320 )  ;
assign n870____DOLLAR__2322 =  ( n510____DOLLAR__1421 ) | ( n869____DOLLAR__2321 )  ;
assign n871____DOLLAR__2323 =  ( n509____DOLLAR__1417 ) | ( n870____DOLLAR__2322 )  ;
assign n872____DOLLAR__2324 =  ( n508____DOLLAR__1413 ) | ( n871____DOLLAR__2323 )  ;
assign n873____DOLLAR__2325 =  ( n507____DOLLAR__1409 ) | ( n872____DOLLAR__2324 )  ;
assign n874____DOLLAR__2326 =  ( n506____DOLLAR__1405 ) | ( n873____DOLLAR__2325 )  ;
assign n875____DOLLAR__2327 =  ( n505____DOLLAR__1401 ) | ( n874____DOLLAR__2326 )  ;
assign n876____DOLLAR__2328 =  ( n504____DOLLAR__1397 ) | ( n875____DOLLAR__2327 )  ;
assign n877____DOLLAR__2329 =  ( n503____DOLLAR__1393 ) | ( n876____DOLLAR__2328 )  ;
assign n878____DOLLAR__2330 =  ( n502____DOLLAR__1389 ) | ( n877____DOLLAR__2329 )  ;
assign n879____DOLLAR__2331 =  ( n501____DOLLAR__1385 ) | ( n878____DOLLAR__2330 )  ;
assign n880____DOLLAR__2332 =  ( n500____DOLLAR__1381 ) | ( n879____DOLLAR__2331 )  ;
assign n881____DOLLAR__2333 =  ( n499____DOLLAR__1377 ) | ( n880____DOLLAR__2332 )  ;
assign n882____DOLLAR__2334 =  ( n498____DOLLAR__1373 ) | ( n881____DOLLAR__2333 )  ;
assign n883____DOLLAR__2335 =  ( n497____DOLLAR__1369 ) | ( n882____DOLLAR__2334 )  ;
assign n884____DOLLAR__2336 =  ( n496____DOLLAR__1365 ) | ( n883____DOLLAR__2335 )  ;
assign n885____DOLLAR__2337 =  ( n495____DOLLAR__1361 ) | ( n884____DOLLAR__2336 )  ;
assign n886____DOLLAR__2338 =  ( n494____DOLLAR__1357 ) | ( n885____DOLLAR__2337 )  ;
assign n887____DOLLAR__2339 =  ( n493____DOLLAR__1353 ) | ( n886____DOLLAR__2338 )  ;
assign n888____DOLLAR__2340 =  ( n492____DOLLAR__1349 ) | ( n887____DOLLAR__2339 )  ;
assign n889____DOLLAR__2341 =  ( n491____DOLLAR__1345 ) | ( n888____DOLLAR__2340 )  ;
assign n890____DOLLAR__2342 =  ( n490____DOLLAR__1341 ) | ( n889____DOLLAR__2341 )  ;
assign n891____DOLLAR__2343 =  ( n489____DOLLAR__1337 ) | ( n890____DOLLAR__2342 )  ;
assign n892____DOLLAR__2344 =  ( n488____DOLLAR__1333 ) | ( n891____DOLLAR__2343 )  ;
assign n893____DOLLAR__2345 =  ( n487____DOLLAR__1329 ) | ( n892____DOLLAR__2344 )  ;
assign n894____DOLLAR__2346 =  ( n486____DOLLAR__1325 ) | ( n893____DOLLAR__2345 )  ;
assign n895____DOLLAR__2347 =  ( n485____DOLLAR__1321 ) | ( n894____DOLLAR__2346 )  ;
assign n896____DOLLAR__2348 =  ( n484____DOLLAR__1317 ) | ( n895____DOLLAR__2347 )  ;
assign n897____DOLLAR__2349 =  ( n483____DOLLAR__1313 ) | ( n896____DOLLAR__2348 )  ;
assign n898____DOLLAR__2350 =  ( n482____DOLLAR__1309 ) | ( n897____DOLLAR__2349 )  ;
assign n899____DOLLAR__2351 =  ( n481____DOLLAR__1305 ) | ( n898____DOLLAR__2350 )  ;
assign n900____DOLLAR__2352 =  ( n480____DOLLAR__1301 ) | ( n899____DOLLAR__2351 )  ;
assign n901____DOLLAR__2353 =  ( n479____DOLLAR__1297 ) | ( n900____DOLLAR__2352 )  ;
assign n902____DOLLAR__2354 =  ( n478____DOLLAR__1293 ) | ( n901____DOLLAR__2353 )  ;
assign n903____DOLLAR__2355 =  ( n477____DOLLAR__1289 ) | ( n902____DOLLAR__2354 )  ;
assign n904____DOLLAR__2356 =  ( n476____DOLLAR__1285 ) | ( n903____DOLLAR__2355 )  ;
assign n905____DOLLAR__2357 =  ( n475____DOLLAR__1281 ) | ( n904____DOLLAR__2356 )  ;
assign n906____DOLLAR__2358 =  ( n474____DOLLAR__1277 ) | ( n905____DOLLAR__2357 )  ;
assign n907____DOLLAR__2359 =  ( n473____DOLLAR__1273 ) | ( n906____DOLLAR__2358 )  ;
assign n908____DOLLAR__2360 =  ( n472____DOLLAR__1269 ) | ( n907____DOLLAR__2359 )  ;
assign n909____DOLLAR__2361 =  ( n471____DOLLAR__1265 ) | ( n908____DOLLAR__2360 )  ;
assign n910____DOLLAR__2362 =  ( n470____DOLLAR__1261 ) | ( n909____DOLLAR__2361 )  ;
assign n911____DOLLAR__2363 =  ( n469____DOLLAR__1257 ) | ( n910____DOLLAR__2362 )  ;
assign n912____DOLLAR__2364 =  ( n468____DOLLAR__1253 ) | ( n911____DOLLAR__2363 )  ;
assign n913____DOLLAR__2365 =  ( n467____DOLLAR__1249 ) | ( n912____DOLLAR__2364 )  ;
assign n914____DOLLAR__2366 =  ( n466____DOLLAR__1245 ) | ( n913____DOLLAR__2365 )  ;
assign n915____DOLLAR__2367 =  ( n465____DOLLAR__1241 ) | ( n914____DOLLAR__2366 )  ;
assign n916____DOLLAR__2368 =  ( n464____DOLLAR__1237 ) | ( n915____DOLLAR__2367 )  ;
assign n917____DOLLAR__2371 = PSW[4:3] ;
assign n918____DOLLAR__2379 =  { ( n917____DOLLAR__2371 ) , ( 3'd7 ) }  ;
assign n919____DOLLAR__2385 =  { ( 3'd0 ) , ( n918____DOLLAR__2379 ) }  ;
assign n920____DOLLAR__2389 =  ( n919____DOLLAR__2385 ) == ( 8'd176 )  ;
assign n921____DOLLAR__2391 =  ( n920____DOLLAR__2389 ) ? ( ACC ) : ( P3 ) ;
assign n922____DOLLAR__2392 =  ( n916____DOLLAR__2368 ) ? ( n921____DOLLAR__2391 ) : ( P3 ) ;
assign n923____DOLLAR__2397 =  ( oc8051_ROM_rdata_0 ) == ( 8'd50 )  ;
assign n924____DOLLAR__2401 =  ( oc8051_ROM_rdata_0 ) == ( 8'd34 )  ;
assign n925____DOLLAR__2403 =  ( n923____DOLLAR__2397 ) | ( n924____DOLLAR__2401 )  ;
assign n926____DOLLAR__177450 = SP[3:0] ;
assign n927____DOLLAR__177531 =  ( n926____DOLLAR__177450 ) == ( 4'd15 )  ;
assign n928____DOLLAR__177526 =  ( n926____DOLLAR__177450 ) == ( 4'd14 )  ;
assign n929____DOLLAR__177521 =  ( n926____DOLLAR__177450 ) == ( 4'd13 )  ;
assign n930____DOLLAR__177516 =  ( n926____DOLLAR__177450 ) == ( 4'd12 )  ;
assign n931____DOLLAR__177511 =  ( n926____DOLLAR__177450 ) == ( 4'd11 )  ;
assign n932____DOLLAR__177506 =  ( n926____DOLLAR__177450 ) == ( 4'd10 )  ;
assign n933____DOLLAR__177501 =  ( n926____DOLLAR__177450 ) == ( 4'd9 )  ;
assign n934____DOLLAR__177496 =  ( n926____DOLLAR__177450 ) == ( 4'd8 )  ;
assign n935____DOLLAR__177491 =  ( n926____DOLLAR__177450 ) == ( 4'd7 )  ;
assign n936____DOLLAR__177486 =  ( n926____DOLLAR__177450 ) == ( 4'd6 )  ;
assign n937____DOLLAR__177481 =  ( n926____DOLLAR__177450 ) == ( 4'd5 )  ;
assign n938____DOLLAR__177476 =  ( n926____DOLLAR__177450 ) == ( 4'd4 )  ;
assign n939____DOLLAR__177471 =  ( n926____DOLLAR__177450 ) == ( 4'd3 )  ;
assign n940____DOLLAR__177466 =  ( n926____DOLLAR__177450 ) == ( 4'd2 )  ;
assign n941____DOLLAR__177461 =  ( n926____DOLLAR__177450 ) == ( 4'd1 )  ;
assign n942____DOLLAR__177456 =  ( n926____DOLLAR__177450 ) == ( 4'd0 )  ;
assign n943____DOLLAR__177458 =  ( n942____DOLLAR__177456 ) ? ( oc8051_IRAM_data_0 ) : ( 8'd0 ) ;
assign n944____DOLLAR__177463 =  ( n941____DOLLAR__177461 ) ? ( oc8051_IRAM_data_1 ) : ( n943____DOLLAR__177458 ) ;
assign n945____DOLLAR__177468 =  ( n940____DOLLAR__177466 ) ? ( oc8051_IRAM_data_2 ) : ( n944____DOLLAR__177463 ) ;
assign n946____DOLLAR__177473 =  ( n939____DOLLAR__177471 ) ? ( oc8051_IRAM_data_3 ) : ( n945____DOLLAR__177468 ) ;
assign n947____DOLLAR__177478 =  ( n938____DOLLAR__177476 ) ? ( oc8051_IRAM_data_4 ) : ( n946____DOLLAR__177473 ) ;
assign n948____DOLLAR__177483 =  ( n937____DOLLAR__177481 ) ? ( oc8051_IRAM_data_5 ) : ( n947____DOLLAR__177478 ) ;
assign n949____DOLLAR__177488 =  ( n936____DOLLAR__177486 ) ? ( oc8051_IRAM_data_6 ) : ( n948____DOLLAR__177483 ) ;
assign n950____DOLLAR__177493 =  ( n935____DOLLAR__177491 ) ? ( oc8051_IRAM_data_7 ) : ( n949____DOLLAR__177488 ) ;
assign n951____DOLLAR__177498 =  ( n934____DOLLAR__177496 ) ? ( oc8051_IRAM_data_8 ) : ( n950____DOLLAR__177493 ) ;
assign n952____DOLLAR__177503 =  ( n933____DOLLAR__177501 ) ? ( oc8051_IRAM_data_9 ) : ( n951____DOLLAR__177498 ) ;
assign n953____DOLLAR__177508 =  ( n932____DOLLAR__177506 ) ? ( oc8051_IRAM_data_10 ) : ( n952____DOLLAR__177503 ) ;
assign n954____DOLLAR__177513 =  ( n931____DOLLAR__177511 ) ? ( oc8051_IRAM_data_11 ) : ( n953____DOLLAR__177508 ) ;
assign n955____DOLLAR__177518 =  ( n930____DOLLAR__177516 ) ? ( oc8051_IRAM_data_12 ) : ( n954____DOLLAR__177513 ) ;
assign n956____DOLLAR__177523 =  ( n929____DOLLAR__177521 ) ? ( oc8051_IRAM_data_13 ) : ( n955____DOLLAR__177518 ) ;
assign n957____DOLLAR__177528 =  ( n928____DOLLAR__177526 ) ? ( oc8051_IRAM_data_14 ) : ( n956____DOLLAR__177523 ) ;
assign n958____DOLLAR__177533 =  ( n927____DOLLAR__177531 ) ? ( oc8051_IRAM_data_15 ) : ( n957____DOLLAR__177528 ) ;
assign n959____DOLLAR__2408 =  ( SP ) - ( 8'd1 )  ;
assign n960____DOLLAR__177535 = n959____DOLLAR__2408[3:0] ;
assign n961____DOLLAR__177616 =  ( n960____DOLLAR__177535 ) == ( 4'd15 )  ;
assign n962____DOLLAR__177611 =  ( n960____DOLLAR__177535 ) == ( 4'd14 )  ;
assign n963____DOLLAR__177606 =  ( n960____DOLLAR__177535 ) == ( 4'd13 )  ;
assign n964____DOLLAR__177601 =  ( n960____DOLLAR__177535 ) == ( 4'd12 )  ;
assign n965____DOLLAR__177596 =  ( n960____DOLLAR__177535 ) == ( 4'd11 )  ;
assign n966____DOLLAR__177591 =  ( n960____DOLLAR__177535 ) == ( 4'd10 )  ;
assign n967____DOLLAR__177586 =  ( n960____DOLLAR__177535 ) == ( 4'd9 )  ;
assign n968____DOLLAR__177581 =  ( n960____DOLLAR__177535 ) == ( 4'd8 )  ;
assign n969____DOLLAR__177576 =  ( n960____DOLLAR__177535 ) == ( 4'd7 )  ;
assign n970____DOLLAR__177571 =  ( n960____DOLLAR__177535 ) == ( 4'd6 )  ;
assign n971____DOLLAR__177566 =  ( n960____DOLLAR__177535 ) == ( 4'd5 )  ;
assign n972____DOLLAR__177561 =  ( n960____DOLLAR__177535 ) == ( 4'd4 )  ;
assign n973____DOLLAR__177556 =  ( n960____DOLLAR__177535 ) == ( 4'd3 )  ;
assign n974____DOLLAR__177551 =  ( n960____DOLLAR__177535 ) == ( 4'd2 )  ;
assign n975____DOLLAR__177546 =  ( n960____DOLLAR__177535 ) == ( 4'd1 )  ;
assign n976____DOLLAR__177541 =  ( n960____DOLLAR__177535 ) == ( 4'd0 )  ;
assign n977____DOLLAR__177543 =  ( n976____DOLLAR__177541 ) ? ( oc8051_IRAM_data_0 ) : ( 8'd0 ) ;
assign n978____DOLLAR__177548 =  ( n975____DOLLAR__177546 ) ? ( oc8051_IRAM_data_1 ) : ( n977____DOLLAR__177543 ) ;
assign n979____DOLLAR__177553 =  ( n974____DOLLAR__177551 ) ? ( oc8051_IRAM_data_2 ) : ( n978____DOLLAR__177548 ) ;
assign n980____DOLLAR__177558 =  ( n973____DOLLAR__177556 ) ? ( oc8051_IRAM_data_3 ) : ( n979____DOLLAR__177553 ) ;
assign n981____DOLLAR__177563 =  ( n972____DOLLAR__177561 ) ? ( oc8051_IRAM_data_4 ) : ( n980____DOLLAR__177558 ) ;
assign n982____DOLLAR__177568 =  ( n971____DOLLAR__177566 ) ? ( oc8051_IRAM_data_5 ) : ( n981____DOLLAR__177563 ) ;
assign n983____DOLLAR__177573 =  ( n970____DOLLAR__177571 ) ? ( oc8051_IRAM_data_6 ) : ( n982____DOLLAR__177568 ) ;
assign n984____DOLLAR__177578 =  ( n969____DOLLAR__177576 ) ? ( oc8051_IRAM_data_7 ) : ( n983____DOLLAR__177573 ) ;
assign n985____DOLLAR__177583 =  ( n968____DOLLAR__177581 ) ? ( oc8051_IRAM_data_8 ) : ( n984____DOLLAR__177578 ) ;
assign n986____DOLLAR__177588 =  ( n967____DOLLAR__177586 ) ? ( oc8051_IRAM_data_9 ) : ( n985____DOLLAR__177583 ) ;
assign n987____DOLLAR__177593 =  ( n966____DOLLAR__177591 ) ? ( oc8051_IRAM_data_10 ) : ( n986____DOLLAR__177588 ) ;
assign n988____DOLLAR__177598 =  ( n965____DOLLAR__177596 ) ? ( oc8051_IRAM_data_11 ) : ( n987____DOLLAR__177593 ) ;
assign n989____DOLLAR__177603 =  ( n964____DOLLAR__177601 ) ? ( oc8051_IRAM_data_12 ) : ( n988____DOLLAR__177598 ) ;
assign n990____DOLLAR__177608 =  ( n963____DOLLAR__177606 ) ? ( oc8051_IRAM_data_13 ) : ( n989____DOLLAR__177603 ) ;
assign n991____DOLLAR__177613 =  ( n962____DOLLAR__177611 ) ? ( oc8051_IRAM_data_14 ) : ( n990____DOLLAR__177608 ) ;
assign n992____DOLLAR__177618 =  ( n961____DOLLAR__177616 ) ? ( oc8051_IRAM_data_15 ) : ( n991____DOLLAR__177613 ) ;
assign n993____DOLLAR__2415 =  { ( n958____DOLLAR__177533 ) , ( n992____DOLLAR__177618 ) }  ;
assign n994____DOLLAR__2421 =  ( oc8051_ROM_rdata_0 ) == ( 8'd49 )  ;
assign n995____DOLLAR__2425 =  ( oc8051_ROM_rdata_0 ) == ( 8'd33 )  ;
assign n996____DOLLAR__2427 =  ( n994____DOLLAR__2421 ) | ( n995____DOLLAR__2425 )  ;
assign n997____DOLLAR__2430 =  ( PC ) + ( 16'd2 )  ;
assign n998____DOLLAR__2431 = n997____DOLLAR__2430[15:11] ;
assign n999____DOLLAR__2439 =  { ( n998____DOLLAR__2431 ) , ( 3'd1 ) }  ;
assign n1000____DOLLAR__2450 =  { ( n999____DOLLAR__2439 ) , ( oc8051_ROM_rdata_1 ) }  ;
assign n1001____DOLLAR__2456 =  ( oc8051_ROM_rdata_0 ) == ( 8'd32 )  ;
assign n1002____DOLLAR__2460 =  ( oc8051_ROM_rdata_0 ) == ( 8'd16 )  ;
assign n1003____DOLLAR__2462 =  ( n1001____DOLLAR__2456 ) | ( n1002____DOLLAR__2460 )  ;
assign n1004____DOLLAR__2468 = oc8051_ROM_rdata_1[7:7] ;
assign n1005____DOLLAR__2472 =  ( n1004____DOLLAR__2468 ) == ( 1'd1 )  ;
assign n1006____DOLLAR__2474 = oc8051_ROM_rdata_1[7:3] ;
assign n1007____DOLLAR__2482 =  { ( n1006____DOLLAR__2474 ) , ( 3'd0 ) }  ;
assign n1008____DOLLAR__2484 =  {3'd0 , n1006____DOLLAR__2474}  ;
assign n1009____DOLLAR__2488 =  ( n1008____DOLLAR__2484 ) + ( 8'd32 )  ;
assign n1010____DOLLAR__2489 =  ( n1005____DOLLAR__2472 ) ? ( n1007____DOLLAR__2482 ) : ( n1009____DOLLAR__2488 ) ;
assign n1011____DOLLAR__2490 = n1010____DOLLAR__2489[7:7] ;
assign n1012____DOLLAR__2494 =  ( n1011____DOLLAR__2490 ) == ( 1'd0 )  ;
assign n1013____DOLLAR__178417 = n1010____DOLLAR__2489[3:0] ;
assign n1014____DOLLAR__178498 =  ( n1013____DOLLAR__178417 ) == ( 4'd15 )  ;
assign n1015____DOLLAR__178493 =  ( n1013____DOLLAR__178417 ) == ( 4'd14 )  ;
assign n1016____DOLLAR__178488 =  ( n1013____DOLLAR__178417 ) == ( 4'd13 )  ;
assign n1017____DOLLAR__178483 =  ( n1013____DOLLAR__178417 ) == ( 4'd12 )  ;
assign n1018____DOLLAR__178478 =  ( n1013____DOLLAR__178417 ) == ( 4'd11 )  ;
assign n1019____DOLLAR__178473 =  ( n1013____DOLLAR__178417 ) == ( 4'd10 )  ;
assign n1020____DOLLAR__178468 =  ( n1013____DOLLAR__178417 ) == ( 4'd9 )  ;
assign n1021____DOLLAR__178463 =  ( n1013____DOLLAR__178417 ) == ( 4'd8 )  ;
assign n1022____DOLLAR__178458 =  ( n1013____DOLLAR__178417 ) == ( 4'd7 )  ;
assign n1023____DOLLAR__178453 =  ( n1013____DOLLAR__178417 ) == ( 4'd6 )  ;
assign n1024____DOLLAR__178448 =  ( n1013____DOLLAR__178417 ) == ( 4'd5 )  ;
assign n1025____DOLLAR__178443 =  ( n1013____DOLLAR__178417 ) == ( 4'd4 )  ;
assign n1026____DOLLAR__178438 =  ( n1013____DOLLAR__178417 ) == ( 4'd3 )  ;
assign n1027____DOLLAR__178433 =  ( n1013____DOLLAR__178417 ) == ( 4'd2 )  ;
assign n1028____DOLLAR__178428 =  ( n1013____DOLLAR__178417 ) == ( 4'd1 )  ;
assign n1029____DOLLAR__178423 =  ( n1013____DOLLAR__178417 ) == ( 4'd0 )  ;
assign n1030____DOLLAR__178425 =  ( n1029____DOLLAR__178423 ) ? ( oc8051_IRAM_data_0 ) : ( 8'd0 ) ;
assign n1031____DOLLAR__178430 =  ( n1028____DOLLAR__178428 ) ? ( oc8051_IRAM_data_1 ) : ( n1030____DOLLAR__178425 ) ;
assign n1032____DOLLAR__178435 =  ( n1027____DOLLAR__178433 ) ? ( oc8051_IRAM_data_2 ) : ( n1031____DOLLAR__178430 ) ;
assign n1033____DOLLAR__178440 =  ( n1026____DOLLAR__178438 ) ? ( oc8051_IRAM_data_3 ) : ( n1032____DOLLAR__178435 ) ;
assign n1034____DOLLAR__178445 =  ( n1025____DOLLAR__178443 ) ? ( oc8051_IRAM_data_4 ) : ( n1033____DOLLAR__178440 ) ;
assign n1035____DOLLAR__178450 =  ( n1024____DOLLAR__178448 ) ? ( oc8051_IRAM_data_5 ) : ( n1034____DOLLAR__178445 ) ;
assign n1036____DOLLAR__178455 =  ( n1023____DOLLAR__178453 ) ? ( oc8051_IRAM_data_6 ) : ( n1035____DOLLAR__178450 ) ;
assign n1037____DOLLAR__178460 =  ( n1022____DOLLAR__178458 ) ? ( oc8051_IRAM_data_7 ) : ( n1036____DOLLAR__178455 ) ;
assign n1038____DOLLAR__178465 =  ( n1021____DOLLAR__178463 ) ? ( oc8051_IRAM_data_8 ) : ( n1037____DOLLAR__178460 ) ;
assign n1039____DOLLAR__178470 =  ( n1020____DOLLAR__178468 ) ? ( oc8051_IRAM_data_9 ) : ( n1038____DOLLAR__178465 ) ;
assign n1040____DOLLAR__178475 =  ( n1019____DOLLAR__178473 ) ? ( oc8051_IRAM_data_10 ) : ( n1039____DOLLAR__178470 ) ;
assign n1041____DOLLAR__178480 =  ( n1018____DOLLAR__178478 ) ? ( oc8051_IRAM_data_11 ) : ( n1040____DOLLAR__178475 ) ;
assign n1042____DOLLAR__178485 =  ( n1017____DOLLAR__178483 ) ? ( oc8051_IRAM_data_12 ) : ( n1041____DOLLAR__178480 ) ;
assign n1043____DOLLAR__178490 =  ( n1016____DOLLAR__178488 ) ? ( oc8051_IRAM_data_13 ) : ( n1042____DOLLAR__178485 ) ;
assign n1044____DOLLAR__178495 =  ( n1015____DOLLAR__178493 ) ? ( oc8051_IRAM_data_14 ) : ( n1043____DOLLAR__178490 ) ;
assign n1045____DOLLAR__178500 =  ( n1014____DOLLAR__178498 ) ? ( oc8051_IRAM_data_15 ) : ( n1044____DOLLAR__178495 ) ;
assign n1046____DOLLAR__2500 =  ( n1010____DOLLAR__2489 ) == ( 8'd128 )  ;
assign n1047____DOLLAR__2504 =  ( n1010____DOLLAR__2489 ) == ( 8'd129 )  ;
assign n1048____DOLLAR__2508 =  ( n1010____DOLLAR__2489 ) == ( 8'd130 )  ;
assign n1049____DOLLAR__2512 =  ( n1010____DOLLAR__2489 ) == ( 8'd131 )  ;
assign n1050____DOLLAR__2516 =  ( n1010____DOLLAR__2489 ) == ( 8'd135 )  ;
assign n1051____DOLLAR__2520 =  ( n1010____DOLLAR__2489 ) == ( 8'd136 )  ;
assign n1052____DOLLAR__2524 =  ( n1010____DOLLAR__2489 ) == ( 8'd137 )  ;
assign n1053____DOLLAR__2528 =  ( n1010____DOLLAR__2489 ) == ( 8'd138 )  ;
assign n1054____DOLLAR__2532 =  ( n1010____DOLLAR__2489 ) == ( 8'd140 )  ;
assign n1055____DOLLAR__2536 =  ( n1010____DOLLAR__2489 ) == ( 8'd139 )  ;
assign n1056____DOLLAR__2540 =  ( n1010____DOLLAR__2489 ) == ( 8'd141 )  ;
assign n1057____DOLLAR__2544 =  ( n1010____DOLLAR__2489 ) == ( 8'd144 )  ;
assign n1058____DOLLAR__2548 =  ( n1010____DOLLAR__2489 ) == ( 8'd152 )  ;
assign n1059____DOLLAR__2552 =  ( n1010____DOLLAR__2489 ) == ( 8'd153 )  ;
assign n1060____DOLLAR__2556 =  ( n1010____DOLLAR__2489 ) == ( 8'd160 )  ;
assign n1061____DOLLAR__2560 =  ( n1010____DOLLAR__2489 ) == ( 8'd168 )  ;
assign n1062____DOLLAR__2564 =  ( n1010____DOLLAR__2489 ) == ( 8'd176 )  ;
assign n1063____DOLLAR__2568 =  ( n1010____DOLLAR__2489 ) == ( 8'd184 )  ;
assign n1064____DOLLAR__2572 =  ( n1010____DOLLAR__2489 ) == ( 8'd208 )  ;
assign n1065____DOLLAR__2576 =  ( n1010____DOLLAR__2489 ) == ( 8'd224 )  ;
assign n1066____DOLLAR__2580 =  ( n1010____DOLLAR__2489 ) == ( 8'd240 )  ;
assign n1067____DOLLAR__2584 =  ( n1066____DOLLAR__2580 ) ? ( B ) : ( 8'd0 ) ;
assign n1068____DOLLAR__2585 =  ( n1065____DOLLAR__2576 ) ? ( ACC ) : ( n1067____DOLLAR__2584 ) ;
assign n1069____DOLLAR__2586 =  ( n1064____DOLLAR__2572 ) ? ( PSW ) : ( n1068____DOLLAR__2585 ) ;
assign n1070____DOLLAR__2587 =  ( n1063____DOLLAR__2568 ) ? ( IP ) : ( n1069____DOLLAR__2586 ) ;
assign n1071____DOLLAR__2588 =  ( n1062____DOLLAR__2564 ) ? ( P3 ) : ( n1070____DOLLAR__2587 ) ;
assign n1072____DOLLAR__2589 =  ( n1061____DOLLAR__2560 ) ? ( IE ) : ( n1071____DOLLAR__2588 ) ;
assign n1073____DOLLAR__2590 =  ( n1060____DOLLAR__2556 ) ? ( P2 ) : ( n1072____DOLLAR__2589 ) ;
assign n1074____DOLLAR__2591 =  ( n1059____DOLLAR__2552 ) ? ( SBUF ) : ( n1073____DOLLAR__2590 ) ;
assign n1075____DOLLAR__2592 =  ( n1058____DOLLAR__2548 ) ? ( SCON ) : ( n1074____DOLLAR__2591 ) ;
assign n1076____DOLLAR__2593 =  ( n1057____DOLLAR__2544 ) ? ( P1 ) : ( n1075____DOLLAR__2592 ) ;
assign n1077____DOLLAR__2594 =  ( n1056____DOLLAR__2540 ) ? ( TH1 ) : ( n1076____DOLLAR__2593 ) ;
assign n1078____DOLLAR__2595 =  ( n1055____DOLLAR__2536 ) ? ( TL1 ) : ( n1077____DOLLAR__2594 ) ;
assign n1079____DOLLAR__2596 =  ( n1054____DOLLAR__2532 ) ? ( TH0 ) : ( n1078____DOLLAR__2595 ) ;
assign n1080____DOLLAR__2597 =  ( n1053____DOLLAR__2528 ) ? ( TL0 ) : ( n1079____DOLLAR__2596 ) ;
assign n1081____DOLLAR__2598 =  ( n1052____DOLLAR__2524 ) ? ( TMOD ) : ( n1080____DOLLAR__2597 ) ;
assign n1082____DOLLAR__2599 =  ( n1051____DOLLAR__2520 ) ? ( TCON ) : ( n1081____DOLLAR__2598 ) ;
assign n1083____DOLLAR__2600 =  ( n1050____DOLLAR__2516 ) ? ( PCON ) : ( n1082____DOLLAR__2599 ) ;
assign n1084____DOLLAR__2601 =  ( n1049____DOLLAR__2512 ) ? ( DPH ) : ( n1083____DOLLAR__2600 ) ;
assign n1085____DOLLAR__2602 =  ( n1048____DOLLAR__2508 ) ? ( DPL ) : ( n1084____DOLLAR__2601 ) ;
assign n1086____DOLLAR__2603 =  ( n1047____DOLLAR__2504 ) ? ( SP ) : ( n1085____DOLLAR__2602 ) ;
assign n1087____DOLLAR__2604 =  ( n1046____DOLLAR__2500 ) ? ( P0 ) : ( n1086____DOLLAR__2603 ) ;
assign n1088____DOLLAR__2605 =  ( n1012____DOLLAR__2494 ) ? ( n1045____DOLLAR__178500 ) : ( n1087____DOLLAR__2604 ) ;
assign n1089____DOLLAR__2606 = n1088____DOLLAR__2605[0:0] ;
assign n1090____DOLLAR__2608 =  ( n1089____DOLLAR__2606 ) == ( 1'd1 )  ;
assign n1091____DOLLAR__2612 =  ( PC ) + ( 16'd3 )  ;
assign n1092____DOLLAR__2618 =  { {8{oc8051_ROM_rdata_2[7] }  }, oc8051_ROM_rdata_2}  ;
assign n1093____DOLLAR__2620 =  ( n1091____DOLLAR__2612 ) + ( n1092____DOLLAR__2618 )  ;
assign n1094____DOLLAR__2623 =  ( PC ) + ( 16'd3 )  ;
assign n1095____DOLLAR__2624 =  ( n1090____DOLLAR__2608 ) ? ( n1093____DOLLAR__2620 ) : ( n1094____DOLLAR__2623 ) ;
assign n1096____DOLLAR__2629 =  ( oc8051_ROM_rdata_0 ) == ( 8'd245 )  ;
assign n1097____DOLLAR__2633 =  ( oc8051_ROM_rdata_0 ) == ( 8'd229 )  ;
assign n1098____DOLLAR__2637 =  ( oc8051_ROM_rdata_0 ) == ( 8'd210 )  ;
assign n1099____DOLLAR__2641 =  ( oc8051_ROM_rdata_0 ) == ( 8'd208 )  ;
assign n1100____DOLLAR__2645 =  ( oc8051_ROM_rdata_0 ) == ( 8'd197 )  ;
assign n1101____DOLLAR__2649 =  ( oc8051_ROM_rdata_0 ) == ( 8'd194 )  ;
assign n1102____DOLLAR__2653 =  ( oc8051_ROM_rdata_0 ) == ( 8'd192 )  ;
assign n1103____DOLLAR__2657 =  ( oc8051_ROM_rdata_0 ) == ( 8'd178 )  ;
assign n1104____DOLLAR__2661 =  ( oc8051_ROM_rdata_0 ) == ( 8'd176 )  ;
assign n1105____DOLLAR__2665 =  ( oc8051_ROM_rdata_0 ) == ( 8'd175 )  ;
assign n1106____DOLLAR__2669 =  ( oc8051_ROM_rdata_0 ) == ( 8'd174 )  ;
assign n1107____DOLLAR__2673 =  ( oc8051_ROM_rdata_0 ) == ( 8'd173 )  ;
assign n1108____DOLLAR__2677 =  ( oc8051_ROM_rdata_0 ) == ( 8'd172 )  ;
assign n1109____DOLLAR__2681 =  ( oc8051_ROM_rdata_0 ) == ( 8'd171 )  ;
assign n1110____DOLLAR__2685 =  ( oc8051_ROM_rdata_0 ) == ( 8'd170 )  ;
assign n1111____DOLLAR__2689 =  ( oc8051_ROM_rdata_0 ) == ( 8'd169 )  ;
assign n1112____DOLLAR__2693 =  ( oc8051_ROM_rdata_0 ) == ( 8'd168 )  ;
assign n1113____DOLLAR__2697 =  ( oc8051_ROM_rdata_0 ) == ( 8'd167 )  ;
assign n1114____DOLLAR__2701 =  ( oc8051_ROM_rdata_0 ) == ( 8'd166 )  ;
assign n1115____DOLLAR__2705 =  ( oc8051_ROM_rdata_0 ) == ( 8'd162 )  ;
assign n1116____DOLLAR__2709 =  ( oc8051_ROM_rdata_0 ) == ( 8'd160 )  ;
assign n1117____DOLLAR__2713 =  ( oc8051_ROM_rdata_0 ) == ( 8'd149 )  ;
assign n1118____DOLLAR__2717 =  ( oc8051_ROM_rdata_0 ) == ( 8'd148 )  ;
assign n1119____DOLLAR__2721 =  ( oc8051_ROM_rdata_0 ) == ( 8'd146 )  ;
assign n1120____DOLLAR__2725 =  ( oc8051_ROM_rdata_0 ) == ( 8'd143 )  ;
assign n1121____DOLLAR__2729 =  ( oc8051_ROM_rdata_0 ) == ( 8'd142 )  ;
assign n1122____DOLLAR__2733 =  ( oc8051_ROM_rdata_0 ) == ( 8'd141 )  ;
assign n1123____DOLLAR__2737 =  ( oc8051_ROM_rdata_0 ) == ( 8'd140 )  ;
assign n1124____DOLLAR__2741 =  ( oc8051_ROM_rdata_0 ) == ( 8'd139 )  ;
assign n1125____DOLLAR__2745 =  ( oc8051_ROM_rdata_0 ) == ( 8'd138 )  ;
assign n1126____DOLLAR__2749 =  ( oc8051_ROM_rdata_0 ) == ( 8'd137 )  ;
assign n1127____DOLLAR__2753 =  ( oc8051_ROM_rdata_0 ) == ( 8'd136 )  ;
assign n1128____DOLLAR__2757 =  ( oc8051_ROM_rdata_0 ) == ( 8'd135 )  ;
assign n1129____DOLLAR__2761 =  ( oc8051_ROM_rdata_0 ) == ( 8'd134 )  ;
assign n1130____DOLLAR__2765 =  ( oc8051_ROM_rdata_0 ) == ( 8'd130 )  ;
assign n1131____DOLLAR__2769 =  ( oc8051_ROM_rdata_0 ) == ( 8'd127 )  ;
assign n1132____DOLLAR__2773 =  ( oc8051_ROM_rdata_0 ) == ( 8'd126 )  ;
assign n1133____DOLLAR__2777 =  ( oc8051_ROM_rdata_0 ) == ( 8'd125 )  ;
assign n1134____DOLLAR__2781 =  ( oc8051_ROM_rdata_0 ) == ( 8'd124 )  ;
assign n1135____DOLLAR__2785 =  ( oc8051_ROM_rdata_0 ) == ( 8'd123 )  ;
assign n1136____DOLLAR__2789 =  ( oc8051_ROM_rdata_0 ) == ( 8'd122 )  ;
assign n1137____DOLLAR__2793 =  ( oc8051_ROM_rdata_0 ) == ( 8'd121 )  ;
assign n1138____DOLLAR__2797 =  ( oc8051_ROM_rdata_0 ) == ( 8'd120 )  ;
assign n1139____DOLLAR__2801 =  ( oc8051_ROM_rdata_0 ) == ( 8'd119 )  ;
assign n1140____DOLLAR__2805 =  ( oc8051_ROM_rdata_0 ) == ( 8'd118 )  ;
assign n1141____DOLLAR__2809 =  ( oc8051_ROM_rdata_0 ) == ( 8'd116 )  ;
assign n1142____DOLLAR__2813 =  ( oc8051_ROM_rdata_0 ) == ( 8'd114 )  ;
assign n1143____DOLLAR__2817 =  ( oc8051_ROM_rdata_0 ) == ( 8'd101 )  ;
assign n1144____DOLLAR__2821 =  ( oc8051_ROM_rdata_0 ) == ( 8'd100 )  ;
assign n1145____DOLLAR__2825 =  ( oc8051_ROM_rdata_0 ) == ( 8'd98 )  ;
assign n1146____DOLLAR__2829 =  ( oc8051_ROM_rdata_0 ) == ( 8'd85 )  ;
assign n1147____DOLLAR__2833 =  ( oc8051_ROM_rdata_0 ) == ( 8'd84 )  ;
assign n1148____DOLLAR__2837 =  ( oc8051_ROM_rdata_0 ) == ( 8'd82 )  ;
assign n1149____DOLLAR__2841 =  ( oc8051_ROM_rdata_0 ) == ( 8'd69 )  ;
assign n1150____DOLLAR__2845 =  ( oc8051_ROM_rdata_0 ) == ( 8'd68 )  ;
assign n1151____DOLLAR__2849 =  ( oc8051_ROM_rdata_0 ) == ( 8'd66 )  ;
assign n1152____DOLLAR__2853 =  ( oc8051_ROM_rdata_0 ) == ( 8'd53 )  ;
assign n1153____DOLLAR__2857 =  ( oc8051_ROM_rdata_0 ) == ( 8'd52 )  ;
assign n1154____DOLLAR__2861 =  ( oc8051_ROM_rdata_0 ) == ( 8'd37 )  ;
assign n1155____DOLLAR__2865 =  ( oc8051_ROM_rdata_0 ) == ( 8'd36 )  ;
assign n1156____DOLLAR__2869 =  ( oc8051_ROM_rdata_0 ) == ( 8'd21 )  ;
assign n1157____DOLLAR__2873 =  ( oc8051_ROM_rdata_0 ) == ( 8'd5 )  ;
assign n1158____DOLLAR__2875 =  ( n1156____DOLLAR__2869 ) | ( n1157____DOLLAR__2873 )  ;
assign n1159____DOLLAR__2876 =  ( n1155____DOLLAR__2865 ) | ( n1158____DOLLAR__2875 )  ;
assign n1160____DOLLAR__2877 =  ( n1154____DOLLAR__2861 ) | ( n1159____DOLLAR__2876 )  ;
assign n1161____DOLLAR__2878 =  ( n1153____DOLLAR__2857 ) | ( n1160____DOLLAR__2877 )  ;
assign n1162____DOLLAR__2879 =  ( n1152____DOLLAR__2853 ) | ( n1161____DOLLAR__2878 )  ;
assign n1163____DOLLAR__2880 =  ( n1151____DOLLAR__2849 ) | ( n1162____DOLLAR__2879 )  ;
assign n1164____DOLLAR__2881 =  ( n1150____DOLLAR__2845 ) | ( n1163____DOLLAR__2880 )  ;
assign n1165____DOLLAR__2882 =  ( n1149____DOLLAR__2841 ) | ( n1164____DOLLAR__2881 )  ;
assign n1166____DOLLAR__2883 =  ( n1148____DOLLAR__2837 ) | ( n1165____DOLLAR__2882 )  ;
assign n1167____DOLLAR__2884 =  ( n1147____DOLLAR__2833 ) | ( n1166____DOLLAR__2883 )  ;
assign n1168____DOLLAR__2885 =  ( n1146____DOLLAR__2829 ) | ( n1167____DOLLAR__2884 )  ;
assign n1169____DOLLAR__2886 =  ( n1145____DOLLAR__2825 ) | ( n1168____DOLLAR__2885 )  ;
assign n1170____DOLLAR__2887 =  ( n1144____DOLLAR__2821 ) | ( n1169____DOLLAR__2886 )  ;
assign n1171____DOLLAR__2888 =  ( n1143____DOLLAR__2817 ) | ( n1170____DOLLAR__2887 )  ;
assign n1172____DOLLAR__2889 =  ( n1142____DOLLAR__2813 ) | ( n1171____DOLLAR__2888 )  ;
assign n1173____DOLLAR__2890 =  ( n1141____DOLLAR__2809 ) | ( n1172____DOLLAR__2889 )  ;
assign n1174____DOLLAR__2891 =  ( n1140____DOLLAR__2805 ) | ( n1173____DOLLAR__2890 )  ;
assign n1175____DOLLAR__2892 =  ( n1139____DOLLAR__2801 ) | ( n1174____DOLLAR__2891 )  ;
assign n1176____DOLLAR__2893 =  ( n1138____DOLLAR__2797 ) | ( n1175____DOLLAR__2892 )  ;
assign n1177____DOLLAR__2894 =  ( n1137____DOLLAR__2793 ) | ( n1176____DOLLAR__2893 )  ;
assign n1178____DOLLAR__2895 =  ( n1136____DOLLAR__2789 ) | ( n1177____DOLLAR__2894 )  ;
assign n1179____DOLLAR__2896 =  ( n1135____DOLLAR__2785 ) | ( n1178____DOLLAR__2895 )  ;
assign n1180____DOLLAR__2897 =  ( n1134____DOLLAR__2781 ) | ( n1179____DOLLAR__2896 )  ;
assign n1181____DOLLAR__2898 =  ( n1133____DOLLAR__2777 ) | ( n1180____DOLLAR__2897 )  ;
assign n1182____DOLLAR__2899 =  ( n1132____DOLLAR__2773 ) | ( n1181____DOLLAR__2898 )  ;
assign n1183____DOLLAR__2900 =  ( n1131____DOLLAR__2769 ) | ( n1182____DOLLAR__2899 )  ;
assign n1184____DOLLAR__2901 =  ( n1130____DOLLAR__2765 ) | ( n1183____DOLLAR__2900 )  ;
assign n1185____DOLLAR__2902 =  ( n1129____DOLLAR__2761 ) | ( n1184____DOLLAR__2901 )  ;
assign n1186____DOLLAR__2903 =  ( n1128____DOLLAR__2757 ) | ( n1185____DOLLAR__2902 )  ;
assign n1187____DOLLAR__2904 =  ( n1127____DOLLAR__2753 ) | ( n1186____DOLLAR__2903 )  ;
assign n1188____DOLLAR__2905 =  ( n1126____DOLLAR__2749 ) | ( n1187____DOLLAR__2904 )  ;
assign n1189____DOLLAR__2906 =  ( n1125____DOLLAR__2745 ) | ( n1188____DOLLAR__2905 )  ;
assign n1190____DOLLAR__2907 =  ( n1124____DOLLAR__2741 ) | ( n1189____DOLLAR__2906 )  ;
assign n1191____DOLLAR__2908 =  ( n1123____DOLLAR__2737 ) | ( n1190____DOLLAR__2907 )  ;
assign n1192____DOLLAR__2909 =  ( n1122____DOLLAR__2733 ) | ( n1191____DOLLAR__2908 )  ;
assign n1193____DOLLAR__2910 =  ( n1121____DOLLAR__2729 ) | ( n1192____DOLLAR__2909 )  ;
assign n1194____DOLLAR__2911 =  ( n1120____DOLLAR__2725 ) | ( n1193____DOLLAR__2910 )  ;
assign n1195____DOLLAR__2912 =  ( n1119____DOLLAR__2721 ) | ( n1194____DOLLAR__2911 )  ;
assign n1196____DOLLAR__2913 =  ( n1118____DOLLAR__2717 ) | ( n1195____DOLLAR__2912 )  ;
assign n1197____DOLLAR__2914 =  ( n1117____DOLLAR__2713 ) | ( n1196____DOLLAR__2913 )  ;
assign n1198____DOLLAR__2915 =  ( n1116____DOLLAR__2709 ) | ( n1197____DOLLAR__2914 )  ;
assign n1199____DOLLAR__2916 =  ( n1115____DOLLAR__2705 ) | ( n1198____DOLLAR__2915 )  ;
assign n1200____DOLLAR__2917 =  ( n1114____DOLLAR__2701 ) | ( n1199____DOLLAR__2916 )  ;
assign n1201____DOLLAR__2918 =  ( n1113____DOLLAR__2697 ) | ( n1200____DOLLAR__2917 )  ;
assign n1202____DOLLAR__2919 =  ( n1112____DOLLAR__2693 ) | ( n1201____DOLLAR__2918 )  ;
assign n1203____DOLLAR__2920 =  ( n1111____DOLLAR__2689 ) | ( n1202____DOLLAR__2919 )  ;
assign n1204____DOLLAR__2921 =  ( n1110____DOLLAR__2685 ) | ( n1203____DOLLAR__2920 )  ;
assign n1205____DOLLAR__2922 =  ( n1109____DOLLAR__2681 ) | ( n1204____DOLLAR__2921 )  ;
assign n1206____DOLLAR__2923 =  ( n1108____DOLLAR__2677 ) | ( n1205____DOLLAR__2922 )  ;
assign n1207____DOLLAR__2924 =  ( n1107____DOLLAR__2673 ) | ( n1206____DOLLAR__2923 )  ;
assign n1208____DOLLAR__2925 =  ( n1106____DOLLAR__2669 ) | ( n1207____DOLLAR__2924 )  ;
assign n1209____DOLLAR__2926 =  ( n1105____DOLLAR__2665 ) | ( n1208____DOLLAR__2925 )  ;
assign n1210____DOLLAR__2927 =  ( n1104____DOLLAR__2661 ) | ( n1209____DOLLAR__2926 )  ;
assign n1211____DOLLAR__2928 =  ( n1103____DOLLAR__2657 ) | ( n1210____DOLLAR__2927 )  ;
assign n1212____DOLLAR__2929 =  ( n1102____DOLLAR__2653 ) | ( n1211____DOLLAR__2928 )  ;
assign n1213____DOLLAR__2930 =  ( n1101____DOLLAR__2649 ) | ( n1212____DOLLAR__2929 )  ;
assign n1214____DOLLAR__2931 =  ( n1100____DOLLAR__2645 ) | ( n1213____DOLLAR__2930 )  ;
assign n1215____DOLLAR__2932 =  ( n1099____DOLLAR__2641 ) | ( n1214____DOLLAR__2931 )  ;
assign n1216____DOLLAR__2933 =  ( n1098____DOLLAR__2637 ) | ( n1215____DOLLAR__2932 )  ;
assign n1217____DOLLAR__2934 =  ( n1097____DOLLAR__2633 ) | ( n1216____DOLLAR__2933 )  ;
assign n1218____DOLLAR__2935 =  ( n1096____DOLLAR__2629 ) | ( n1217____DOLLAR__2934 )  ;
assign n1219____DOLLAR__2938 =  ( PC ) + ( 16'd2 )  ;
assign n1220____DOLLAR__2943 =  ( oc8051_ROM_rdata_0 ) == ( 8'd18 )  ;
assign n1221____DOLLAR__2947 =  ( oc8051_ROM_rdata_0 ) == ( 8'd2 )  ;
assign n1222____DOLLAR__2949 =  ( n1220____DOLLAR__2943 ) | ( n1221____DOLLAR__2947 )  ;
assign n1223____DOLLAR__2964 =  { ( oc8051_ROM_rdata_1 ) , ( oc8051_ROM_rdata_2 ) }  ;
assign n1224____DOLLAR__2970 =  ( oc8051_ROM_rdata_0 ) == ( 8'd17 )  ;
assign n1225____DOLLAR__2974 =  ( oc8051_ROM_rdata_0 ) == ( 8'd1 )  ;
assign n1226____DOLLAR__2976 =  ( n1224____DOLLAR__2970 ) | ( n1225____DOLLAR__2974 )  ;
assign n1227____DOLLAR__2979 =  ( PC ) + ( 16'd2 )  ;
assign n1228____DOLLAR__2980 = n1227____DOLLAR__2979[15:11] ;
assign n1229____DOLLAR__2988 =  { ( n1228____DOLLAR__2980 ) , ( 3'd0 ) }  ;
assign n1230____DOLLAR__2999 =  { ( n1229____DOLLAR__2988 ) , ( oc8051_ROM_rdata_1 ) }  ;
assign n1231____DOLLAR__3005 =  ( oc8051_ROM_rdata_0 ) == ( 8'd255 )  ;
assign n1232____DOLLAR__3009 =  ( oc8051_ROM_rdata_0 ) == ( 8'd254 )  ;
assign n1233____DOLLAR__3013 =  ( oc8051_ROM_rdata_0 ) == ( 8'd253 )  ;
assign n1234____DOLLAR__3017 =  ( oc8051_ROM_rdata_0 ) == ( 8'd252 )  ;
assign n1235____DOLLAR__3021 =  ( oc8051_ROM_rdata_0 ) == ( 8'd251 )  ;
assign n1236____DOLLAR__3025 =  ( oc8051_ROM_rdata_0 ) == ( 8'd250 )  ;
assign n1237____DOLLAR__3029 =  ( oc8051_ROM_rdata_0 ) == ( 8'd249 )  ;
assign n1238____DOLLAR__3033 =  ( oc8051_ROM_rdata_0 ) == ( 8'd248 )  ;
assign n1239____DOLLAR__3037 =  ( oc8051_ROM_rdata_0 ) == ( 8'd247 )  ;
assign n1240____DOLLAR__3041 =  ( oc8051_ROM_rdata_0 ) == ( 8'd246 )  ;
assign n1241____DOLLAR__3045 =  ( oc8051_ROM_rdata_0 ) == ( 8'd244 )  ;
assign n1242____DOLLAR__3049 =  ( oc8051_ROM_rdata_0 ) == ( 8'd243 )  ;
assign n1243____DOLLAR__3053 =  ( oc8051_ROM_rdata_0 ) == ( 8'd242 )  ;
assign n1244____DOLLAR__3057 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign n1245____DOLLAR__3061 =  ( oc8051_ROM_rdata_0 ) == ( 8'd239 )  ;
assign n1246____DOLLAR__3065 =  ( oc8051_ROM_rdata_0 ) == ( 8'd238 )  ;
assign n1247____DOLLAR__3069 =  ( oc8051_ROM_rdata_0 ) == ( 8'd237 )  ;
assign n1248____DOLLAR__3073 =  ( oc8051_ROM_rdata_0 ) == ( 8'd236 )  ;
assign n1249____DOLLAR__3077 =  ( oc8051_ROM_rdata_0 ) == ( 8'd235 )  ;
assign n1250____DOLLAR__3081 =  ( oc8051_ROM_rdata_0 ) == ( 8'd234 )  ;
assign n1251____DOLLAR__3085 =  ( oc8051_ROM_rdata_0 ) == ( 8'd233 )  ;
assign n1252____DOLLAR__3089 =  ( oc8051_ROM_rdata_0 ) == ( 8'd232 )  ;
assign n1253____DOLLAR__3093 =  ( oc8051_ROM_rdata_0 ) == ( 8'd231 )  ;
assign n1254____DOLLAR__3097 =  ( oc8051_ROM_rdata_0 ) == ( 8'd230 )  ;
assign n1255____DOLLAR__3101 =  ( oc8051_ROM_rdata_0 ) == ( 8'd228 )  ;
assign n1256____DOLLAR__3105 =  ( oc8051_ROM_rdata_0 ) == ( 8'd227 )  ;
assign n1257____DOLLAR__3109 =  ( oc8051_ROM_rdata_0 ) == ( 8'd226 )  ;
assign n1258____DOLLAR__3113 =  ( oc8051_ROM_rdata_0 ) == ( 8'd224 )  ;
assign n1259____DOLLAR__3117 =  ( oc8051_ROM_rdata_0 ) == ( 8'd215 )  ;
assign n1260____DOLLAR__3121 =  ( oc8051_ROM_rdata_0 ) == ( 8'd214 )  ;
assign n1261____DOLLAR__3125 =  ( oc8051_ROM_rdata_0 ) == ( 8'd212 )  ;
assign n1262____DOLLAR__3129 =  ( oc8051_ROM_rdata_0 ) == ( 8'd211 )  ;
assign n1263____DOLLAR__3133 =  ( oc8051_ROM_rdata_0 ) == ( 8'd207 )  ;
assign n1264____DOLLAR__3137 =  ( oc8051_ROM_rdata_0 ) == ( 8'd206 )  ;
assign n1265____DOLLAR__3141 =  ( oc8051_ROM_rdata_0 ) == ( 8'd205 )  ;
assign n1266____DOLLAR__3145 =  ( oc8051_ROM_rdata_0 ) == ( 8'd204 )  ;
assign n1267____DOLLAR__3149 =  ( oc8051_ROM_rdata_0 ) == ( 8'd203 )  ;
assign n1268____DOLLAR__3153 =  ( oc8051_ROM_rdata_0 ) == ( 8'd202 )  ;
assign n1269____DOLLAR__3157 =  ( oc8051_ROM_rdata_0 ) == ( 8'd201 )  ;
assign n1270____DOLLAR__3161 =  ( oc8051_ROM_rdata_0 ) == ( 8'd200 )  ;
assign n1271____DOLLAR__3165 =  ( oc8051_ROM_rdata_0 ) == ( 8'd199 )  ;
assign n1272____DOLLAR__3169 =  ( oc8051_ROM_rdata_0 ) == ( 8'd198 )  ;
assign n1273____DOLLAR__3173 =  ( oc8051_ROM_rdata_0 ) == ( 8'd196 )  ;
assign n1274____DOLLAR__3177 =  ( oc8051_ROM_rdata_0 ) == ( 8'd195 )  ;
assign n1275____DOLLAR__3181 =  ( oc8051_ROM_rdata_0 ) == ( 8'd179 )  ;
assign n1276____DOLLAR__3185 =  ( oc8051_ROM_rdata_0 ) == ( 8'd165 )  ;
assign n1277____DOLLAR__3189 =  ( oc8051_ROM_rdata_0 ) == ( 8'd164 )  ;
assign n1278____DOLLAR__3193 =  ( oc8051_ROM_rdata_0 ) == ( 8'd163 )  ;
assign n1279____DOLLAR__3197 =  ( oc8051_ROM_rdata_0 ) == ( 8'd159 )  ;
assign n1280____DOLLAR__3201 =  ( oc8051_ROM_rdata_0 ) == ( 8'd158 )  ;
assign n1281____DOLLAR__3205 =  ( oc8051_ROM_rdata_0 ) == ( 8'd157 )  ;
assign n1282____DOLLAR__3209 =  ( oc8051_ROM_rdata_0 ) == ( 8'd156 )  ;
assign n1283____DOLLAR__3213 =  ( oc8051_ROM_rdata_0 ) == ( 8'd155 )  ;
assign n1284____DOLLAR__3217 =  ( oc8051_ROM_rdata_0 ) == ( 8'd154 )  ;
assign n1285____DOLLAR__3221 =  ( oc8051_ROM_rdata_0 ) == ( 8'd153 )  ;
assign n1286____DOLLAR__3225 =  ( oc8051_ROM_rdata_0 ) == ( 8'd152 )  ;
assign n1287____DOLLAR__3229 =  ( oc8051_ROM_rdata_0 ) == ( 8'd151 )  ;
assign n1288____DOLLAR__3233 =  ( oc8051_ROM_rdata_0 ) == ( 8'd150 )  ;
assign n1289____DOLLAR__3237 =  ( oc8051_ROM_rdata_0 ) == ( 8'd147 )  ;
assign n1290____DOLLAR__3241 =  ( oc8051_ROM_rdata_0 ) == ( 8'd132 )  ;
assign n1291____DOLLAR__3245 =  ( oc8051_ROM_rdata_0 ) == ( 8'd131 )  ;
assign n1292____DOLLAR__3249 =  ( oc8051_ROM_rdata_0 ) == ( 8'd111 )  ;
assign n1293____DOLLAR__3253 =  ( oc8051_ROM_rdata_0 ) == ( 8'd110 )  ;
assign n1294____DOLLAR__3257 =  ( oc8051_ROM_rdata_0 ) == ( 8'd109 )  ;
assign n1295____DOLLAR__3261 =  ( oc8051_ROM_rdata_0 ) == ( 8'd108 )  ;
assign n1296____DOLLAR__3265 =  ( oc8051_ROM_rdata_0 ) == ( 8'd107 )  ;
assign n1297____DOLLAR__3269 =  ( oc8051_ROM_rdata_0 ) == ( 8'd106 )  ;
assign n1298____DOLLAR__3273 =  ( oc8051_ROM_rdata_0 ) == ( 8'd105 )  ;
assign n1299____DOLLAR__3277 =  ( oc8051_ROM_rdata_0 ) == ( 8'd104 )  ;
assign n1300____DOLLAR__3281 =  ( oc8051_ROM_rdata_0 ) == ( 8'd103 )  ;
assign n1301____DOLLAR__3285 =  ( oc8051_ROM_rdata_0 ) == ( 8'd102 )  ;
assign n1302____DOLLAR__3289 =  ( oc8051_ROM_rdata_0 ) == ( 8'd95 )  ;
assign n1303____DOLLAR__3293 =  ( oc8051_ROM_rdata_0 ) == ( 8'd94 )  ;
assign n1304____DOLLAR__3297 =  ( oc8051_ROM_rdata_0 ) == ( 8'd93 )  ;
assign n1305____DOLLAR__3301 =  ( oc8051_ROM_rdata_0 ) == ( 8'd92 )  ;
assign n1306____DOLLAR__3305 =  ( oc8051_ROM_rdata_0 ) == ( 8'd91 )  ;
assign n1307____DOLLAR__3309 =  ( oc8051_ROM_rdata_0 ) == ( 8'd90 )  ;
assign n1308____DOLLAR__3313 =  ( oc8051_ROM_rdata_0 ) == ( 8'd89 )  ;
assign n1309____DOLLAR__3317 =  ( oc8051_ROM_rdata_0 ) == ( 8'd88 )  ;
assign n1310____DOLLAR__3321 =  ( oc8051_ROM_rdata_0 ) == ( 8'd87 )  ;
assign n1311____DOLLAR__3325 =  ( oc8051_ROM_rdata_0 ) == ( 8'd86 )  ;
assign n1312____DOLLAR__3329 =  ( oc8051_ROM_rdata_0 ) == ( 8'd79 )  ;
assign n1313____DOLLAR__3333 =  ( oc8051_ROM_rdata_0 ) == ( 8'd78 )  ;
assign n1314____DOLLAR__3337 =  ( oc8051_ROM_rdata_0 ) == ( 8'd77 )  ;
assign n1315____DOLLAR__3341 =  ( oc8051_ROM_rdata_0 ) == ( 8'd76 )  ;
assign n1316____DOLLAR__3345 =  ( oc8051_ROM_rdata_0 ) == ( 8'd75 )  ;
assign n1317____DOLLAR__3349 =  ( oc8051_ROM_rdata_0 ) == ( 8'd74 )  ;
assign n1318____DOLLAR__3353 =  ( oc8051_ROM_rdata_0 ) == ( 8'd73 )  ;
assign n1319____DOLLAR__3357 =  ( oc8051_ROM_rdata_0 ) == ( 8'd72 )  ;
assign n1320____DOLLAR__3361 =  ( oc8051_ROM_rdata_0 ) == ( 8'd71 )  ;
assign n1321____DOLLAR__3365 =  ( oc8051_ROM_rdata_0 ) == ( 8'd70 )  ;
assign n1322____DOLLAR__3369 =  ( oc8051_ROM_rdata_0 ) == ( 8'd63 )  ;
assign n1323____DOLLAR__3373 =  ( oc8051_ROM_rdata_0 ) == ( 8'd62 )  ;
assign n1324____DOLLAR__3377 =  ( oc8051_ROM_rdata_0 ) == ( 8'd61 )  ;
assign n1325____DOLLAR__3381 =  ( oc8051_ROM_rdata_0 ) == ( 8'd60 )  ;
assign n1326____DOLLAR__3385 =  ( oc8051_ROM_rdata_0 ) == ( 8'd59 )  ;
assign n1327____DOLLAR__3389 =  ( oc8051_ROM_rdata_0 ) == ( 8'd58 )  ;
assign n1328____DOLLAR__3393 =  ( oc8051_ROM_rdata_0 ) == ( 8'd57 )  ;
assign n1329____DOLLAR__3397 =  ( oc8051_ROM_rdata_0 ) == ( 8'd56 )  ;
assign n1330____DOLLAR__3401 =  ( oc8051_ROM_rdata_0 ) == ( 8'd55 )  ;
assign n1331____DOLLAR__3405 =  ( oc8051_ROM_rdata_0 ) == ( 8'd54 )  ;
assign n1332____DOLLAR__3409 =  ( oc8051_ROM_rdata_0 ) == ( 8'd51 )  ;
assign n1333____DOLLAR__3413 =  ( oc8051_ROM_rdata_0 ) == ( 8'd47 )  ;
assign n1334____DOLLAR__3417 =  ( oc8051_ROM_rdata_0 ) == ( 8'd46 )  ;
assign n1335____DOLLAR__3421 =  ( oc8051_ROM_rdata_0 ) == ( 8'd45 )  ;
assign n1336____DOLLAR__3425 =  ( oc8051_ROM_rdata_0 ) == ( 8'd44 )  ;
assign n1337____DOLLAR__3429 =  ( oc8051_ROM_rdata_0 ) == ( 8'd43 )  ;
assign n1338____DOLLAR__3433 =  ( oc8051_ROM_rdata_0 ) == ( 8'd42 )  ;
assign n1339____DOLLAR__3437 =  ( oc8051_ROM_rdata_0 ) == ( 8'd41 )  ;
assign n1340____DOLLAR__3441 =  ( oc8051_ROM_rdata_0 ) == ( 8'd40 )  ;
assign n1341____DOLLAR__3445 =  ( oc8051_ROM_rdata_0 ) == ( 8'd39 )  ;
assign n1342____DOLLAR__3449 =  ( oc8051_ROM_rdata_0 ) == ( 8'd38 )  ;
assign n1343____DOLLAR__3453 =  ( oc8051_ROM_rdata_0 ) == ( 8'd35 )  ;
assign n1344____DOLLAR__3457 =  ( oc8051_ROM_rdata_0 ) == ( 8'd31 )  ;
assign n1345____DOLLAR__3461 =  ( oc8051_ROM_rdata_0 ) == ( 8'd30 )  ;
assign n1346____DOLLAR__3465 =  ( oc8051_ROM_rdata_0 ) == ( 8'd29 )  ;
assign n1347____DOLLAR__3469 =  ( oc8051_ROM_rdata_0 ) == ( 8'd28 )  ;
assign n1348____DOLLAR__3473 =  ( oc8051_ROM_rdata_0 ) == ( 8'd27 )  ;
assign n1349____DOLLAR__3477 =  ( oc8051_ROM_rdata_0 ) == ( 8'd26 )  ;
assign n1350____DOLLAR__3481 =  ( oc8051_ROM_rdata_0 ) == ( 8'd25 )  ;
assign n1351____DOLLAR__3485 =  ( oc8051_ROM_rdata_0 ) == ( 8'd24 )  ;
assign n1352____DOLLAR__3489 =  ( oc8051_ROM_rdata_0 ) == ( 8'd23 )  ;
assign n1353____DOLLAR__3493 =  ( oc8051_ROM_rdata_0 ) == ( 8'd22 )  ;
assign n1354____DOLLAR__3497 =  ( oc8051_ROM_rdata_0 ) == ( 8'd20 )  ;
assign n1355____DOLLAR__3501 =  ( oc8051_ROM_rdata_0 ) == ( 8'd19 )  ;
assign n1356____DOLLAR__3505 =  ( oc8051_ROM_rdata_0 ) == ( 8'd15 )  ;
assign n1357____DOLLAR__3509 =  ( oc8051_ROM_rdata_0 ) == ( 8'd14 )  ;
assign n1358____DOLLAR__3513 =  ( oc8051_ROM_rdata_0 ) == ( 8'd13 )  ;
assign n1359____DOLLAR__3517 =  ( oc8051_ROM_rdata_0 ) == ( 8'd12 )  ;
assign n1360____DOLLAR__3521 =  ( oc8051_ROM_rdata_0 ) == ( 8'd11 )  ;
assign n1361____DOLLAR__3525 =  ( oc8051_ROM_rdata_0 ) == ( 8'd10 )  ;
assign n1362____DOLLAR__3529 =  ( oc8051_ROM_rdata_0 ) == ( 8'd9 )  ;
assign n1363____DOLLAR__3533 =  ( oc8051_ROM_rdata_0 ) == ( 8'd8 )  ;
assign n1364____DOLLAR__3537 =  ( oc8051_ROM_rdata_0 ) == ( 8'd7 )  ;
assign n1365____DOLLAR__3541 =  ( oc8051_ROM_rdata_0 ) == ( 8'd6 )  ;
assign n1366____DOLLAR__3545 =  ( oc8051_ROM_rdata_0 ) == ( 8'd4 )  ;
assign n1367____DOLLAR__3549 =  ( oc8051_ROM_rdata_0 ) == ( 8'd3 )  ;
assign n1368____DOLLAR__3553 =  ( oc8051_ROM_rdata_0 ) == ( 8'd0 )  ;
assign n1369____DOLLAR__3555 =  ( n1367____DOLLAR__3549 ) | ( n1368____DOLLAR__3553 )  ;
assign n1370____DOLLAR__3556 =  ( n1366____DOLLAR__3545 ) | ( n1369____DOLLAR__3555 )  ;
assign n1371____DOLLAR__3557 =  ( n1365____DOLLAR__3541 ) | ( n1370____DOLLAR__3556 )  ;
assign n1372____DOLLAR__3558 =  ( n1364____DOLLAR__3537 ) | ( n1371____DOLLAR__3557 )  ;
assign n1373____DOLLAR__3559 =  ( n1363____DOLLAR__3533 ) | ( n1372____DOLLAR__3558 )  ;
assign n1374____DOLLAR__3560 =  ( n1362____DOLLAR__3529 ) | ( n1373____DOLLAR__3559 )  ;
assign n1375____DOLLAR__3561 =  ( n1361____DOLLAR__3525 ) | ( n1374____DOLLAR__3560 )  ;
assign n1376____DOLLAR__3562 =  ( n1360____DOLLAR__3521 ) | ( n1375____DOLLAR__3561 )  ;
assign n1377____DOLLAR__3563 =  ( n1359____DOLLAR__3517 ) | ( n1376____DOLLAR__3562 )  ;
assign n1378____DOLLAR__3564 =  ( n1358____DOLLAR__3513 ) | ( n1377____DOLLAR__3563 )  ;
assign n1379____DOLLAR__3565 =  ( n1357____DOLLAR__3509 ) | ( n1378____DOLLAR__3564 )  ;
assign n1380____DOLLAR__3566 =  ( n1356____DOLLAR__3505 ) | ( n1379____DOLLAR__3565 )  ;
assign n1381____DOLLAR__3567 =  ( n1355____DOLLAR__3501 ) | ( n1380____DOLLAR__3566 )  ;
assign n1382____DOLLAR__3568 =  ( n1354____DOLLAR__3497 ) | ( n1381____DOLLAR__3567 )  ;
assign n1383____DOLLAR__3569 =  ( n1353____DOLLAR__3493 ) | ( n1382____DOLLAR__3568 )  ;
assign n1384____DOLLAR__3570 =  ( n1352____DOLLAR__3489 ) | ( n1383____DOLLAR__3569 )  ;
assign n1385____DOLLAR__3571 =  ( n1351____DOLLAR__3485 ) | ( n1384____DOLLAR__3570 )  ;
assign n1386____DOLLAR__3572 =  ( n1350____DOLLAR__3481 ) | ( n1385____DOLLAR__3571 )  ;
assign n1387____DOLLAR__3573 =  ( n1349____DOLLAR__3477 ) | ( n1386____DOLLAR__3572 )  ;
assign n1388____DOLLAR__3574 =  ( n1348____DOLLAR__3473 ) | ( n1387____DOLLAR__3573 )  ;
assign n1389____DOLLAR__3575 =  ( n1347____DOLLAR__3469 ) | ( n1388____DOLLAR__3574 )  ;
assign n1390____DOLLAR__3576 =  ( n1346____DOLLAR__3465 ) | ( n1389____DOLLAR__3575 )  ;
assign n1391____DOLLAR__3577 =  ( n1345____DOLLAR__3461 ) | ( n1390____DOLLAR__3576 )  ;
assign n1392____DOLLAR__3578 =  ( n1344____DOLLAR__3457 ) | ( n1391____DOLLAR__3577 )  ;
assign n1393____DOLLAR__3579 =  ( n1343____DOLLAR__3453 ) | ( n1392____DOLLAR__3578 )  ;
assign n1394____DOLLAR__3580 =  ( n1342____DOLLAR__3449 ) | ( n1393____DOLLAR__3579 )  ;
assign n1395____DOLLAR__3581 =  ( n1341____DOLLAR__3445 ) | ( n1394____DOLLAR__3580 )  ;
assign n1396____DOLLAR__3582 =  ( n1340____DOLLAR__3441 ) | ( n1395____DOLLAR__3581 )  ;
assign n1397____DOLLAR__3583 =  ( n1339____DOLLAR__3437 ) | ( n1396____DOLLAR__3582 )  ;
assign n1398____DOLLAR__3584 =  ( n1338____DOLLAR__3433 ) | ( n1397____DOLLAR__3583 )  ;
assign n1399____DOLLAR__3585 =  ( n1337____DOLLAR__3429 ) | ( n1398____DOLLAR__3584 )  ;
assign n1400____DOLLAR__3586 =  ( n1336____DOLLAR__3425 ) | ( n1399____DOLLAR__3585 )  ;
assign n1401____DOLLAR__3587 =  ( n1335____DOLLAR__3421 ) | ( n1400____DOLLAR__3586 )  ;
assign n1402____DOLLAR__3588 =  ( n1334____DOLLAR__3417 ) | ( n1401____DOLLAR__3587 )  ;
assign n1403____DOLLAR__3589 =  ( n1333____DOLLAR__3413 ) | ( n1402____DOLLAR__3588 )  ;
assign n1404____DOLLAR__3590 =  ( n1332____DOLLAR__3409 ) | ( n1403____DOLLAR__3589 )  ;
assign n1405____DOLLAR__3591 =  ( n1331____DOLLAR__3405 ) | ( n1404____DOLLAR__3590 )  ;
assign n1406____DOLLAR__3592 =  ( n1330____DOLLAR__3401 ) | ( n1405____DOLLAR__3591 )  ;
assign n1407____DOLLAR__3593 =  ( n1329____DOLLAR__3397 ) | ( n1406____DOLLAR__3592 )  ;
assign n1408____DOLLAR__3594 =  ( n1328____DOLLAR__3393 ) | ( n1407____DOLLAR__3593 )  ;
assign n1409____DOLLAR__3595 =  ( n1327____DOLLAR__3389 ) | ( n1408____DOLLAR__3594 )  ;
assign n1410____DOLLAR__3596 =  ( n1326____DOLLAR__3385 ) | ( n1409____DOLLAR__3595 )  ;
assign n1411____DOLLAR__3597 =  ( n1325____DOLLAR__3381 ) | ( n1410____DOLLAR__3596 )  ;
assign n1412____DOLLAR__3598 =  ( n1324____DOLLAR__3377 ) | ( n1411____DOLLAR__3597 )  ;
assign n1413____DOLLAR__3599 =  ( n1323____DOLLAR__3373 ) | ( n1412____DOLLAR__3598 )  ;
assign n1414____DOLLAR__3600 =  ( n1322____DOLLAR__3369 ) | ( n1413____DOLLAR__3599 )  ;
assign n1415____DOLLAR__3601 =  ( n1321____DOLLAR__3365 ) | ( n1414____DOLLAR__3600 )  ;
assign n1416____DOLLAR__3602 =  ( n1320____DOLLAR__3361 ) | ( n1415____DOLLAR__3601 )  ;
assign n1417____DOLLAR__3603 =  ( n1319____DOLLAR__3357 ) | ( n1416____DOLLAR__3602 )  ;
assign n1418____DOLLAR__3604 =  ( n1318____DOLLAR__3353 ) | ( n1417____DOLLAR__3603 )  ;
assign n1419____DOLLAR__3605 =  ( n1317____DOLLAR__3349 ) | ( n1418____DOLLAR__3604 )  ;
assign n1420____DOLLAR__3606 =  ( n1316____DOLLAR__3345 ) | ( n1419____DOLLAR__3605 )  ;
assign n1421____DOLLAR__3607 =  ( n1315____DOLLAR__3341 ) | ( n1420____DOLLAR__3606 )  ;
assign n1422____DOLLAR__3608 =  ( n1314____DOLLAR__3337 ) | ( n1421____DOLLAR__3607 )  ;
assign n1423____DOLLAR__3609 =  ( n1313____DOLLAR__3333 ) | ( n1422____DOLLAR__3608 )  ;
assign n1424____DOLLAR__3610 =  ( n1312____DOLLAR__3329 ) | ( n1423____DOLLAR__3609 )  ;
assign n1425____DOLLAR__3611 =  ( n1311____DOLLAR__3325 ) | ( n1424____DOLLAR__3610 )  ;
assign n1426____DOLLAR__3612 =  ( n1310____DOLLAR__3321 ) | ( n1425____DOLLAR__3611 )  ;
assign n1427____DOLLAR__3613 =  ( n1309____DOLLAR__3317 ) | ( n1426____DOLLAR__3612 )  ;
assign n1428____DOLLAR__3614 =  ( n1308____DOLLAR__3313 ) | ( n1427____DOLLAR__3613 )  ;
assign n1429____DOLLAR__3615 =  ( n1307____DOLLAR__3309 ) | ( n1428____DOLLAR__3614 )  ;
assign n1430____DOLLAR__3616 =  ( n1306____DOLLAR__3305 ) | ( n1429____DOLLAR__3615 )  ;
assign n1431____DOLLAR__3617 =  ( n1305____DOLLAR__3301 ) | ( n1430____DOLLAR__3616 )  ;
assign n1432____DOLLAR__3618 =  ( n1304____DOLLAR__3297 ) | ( n1431____DOLLAR__3617 )  ;
assign n1433____DOLLAR__3619 =  ( n1303____DOLLAR__3293 ) | ( n1432____DOLLAR__3618 )  ;
assign n1434____DOLLAR__3620 =  ( n1302____DOLLAR__3289 ) | ( n1433____DOLLAR__3619 )  ;
assign n1435____DOLLAR__3621 =  ( n1301____DOLLAR__3285 ) | ( n1434____DOLLAR__3620 )  ;
assign n1436____DOLLAR__3622 =  ( n1300____DOLLAR__3281 ) | ( n1435____DOLLAR__3621 )  ;
assign n1437____DOLLAR__3623 =  ( n1299____DOLLAR__3277 ) | ( n1436____DOLLAR__3622 )  ;
assign n1438____DOLLAR__3624 =  ( n1298____DOLLAR__3273 ) | ( n1437____DOLLAR__3623 )  ;
assign n1439____DOLLAR__3625 =  ( n1297____DOLLAR__3269 ) | ( n1438____DOLLAR__3624 )  ;
assign n1440____DOLLAR__3626 =  ( n1296____DOLLAR__3265 ) | ( n1439____DOLLAR__3625 )  ;
assign n1441____DOLLAR__3627 =  ( n1295____DOLLAR__3261 ) | ( n1440____DOLLAR__3626 )  ;
assign n1442____DOLLAR__3628 =  ( n1294____DOLLAR__3257 ) | ( n1441____DOLLAR__3627 )  ;
assign n1443____DOLLAR__3629 =  ( n1293____DOLLAR__3253 ) | ( n1442____DOLLAR__3628 )  ;
assign n1444____DOLLAR__3630 =  ( n1292____DOLLAR__3249 ) | ( n1443____DOLLAR__3629 )  ;
assign n1445____DOLLAR__3631 =  ( n1291____DOLLAR__3245 ) | ( n1444____DOLLAR__3630 )  ;
assign n1446____DOLLAR__3632 =  ( n1290____DOLLAR__3241 ) | ( n1445____DOLLAR__3631 )  ;
assign n1447____DOLLAR__3633 =  ( n1289____DOLLAR__3237 ) | ( n1446____DOLLAR__3632 )  ;
assign n1448____DOLLAR__3634 =  ( n1288____DOLLAR__3233 ) | ( n1447____DOLLAR__3633 )  ;
assign n1449____DOLLAR__3635 =  ( n1287____DOLLAR__3229 ) | ( n1448____DOLLAR__3634 )  ;
assign n1450____DOLLAR__3636 =  ( n1286____DOLLAR__3225 ) | ( n1449____DOLLAR__3635 )  ;
assign n1451____DOLLAR__3637 =  ( n1285____DOLLAR__3221 ) | ( n1450____DOLLAR__3636 )  ;
assign n1452____DOLLAR__3638 =  ( n1284____DOLLAR__3217 ) | ( n1451____DOLLAR__3637 )  ;
assign n1453____DOLLAR__3639 =  ( n1283____DOLLAR__3213 ) | ( n1452____DOLLAR__3638 )  ;
assign n1454____DOLLAR__3640 =  ( n1282____DOLLAR__3209 ) | ( n1453____DOLLAR__3639 )  ;
assign n1455____DOLLAR__3641 =  ( n1281____DOLLAR__3205 ) | ( n1454____DOLLAR__3640 )  ;
assign n1456____DOLLAR__3642 =  ( n1280____DOLLAR__3201 ) | ( n1455____DOLLAR__3641 )  ;
assign n1457____DOLLAR__3643 =  ( n1279____DOLLAR__3197 ) | ( n1456____DOLLAR__3642 )  ;
assign n1458____DOLLAR__3644 =  ( n1278____DOLLAR__3193 ) | ( n1457____DOLLAR__3643 )  ;
assign n1459____DOLLAR__3645 =  ( n1277____DOLLAR__3189 ) | ( n1458____DOLLAR__3644 )  ;
assign n1460____DOLLAR__3646 =  ( n1276____DOLLAR__3185 ) | ( n1459____DOLLAR__3645 )  ;
assign n1461____DOLLAR__3647 =  ( n1275____DOLLAR__3181 ) | ( n1460____DOLLAR__3646 )  ;
assign n1462____DOLLAR__3648 =  ( n1274____DOLLAR__3177 ) | ( n1461____DOLLAR__3647 )  ;
assign n1463____DOLLAR__3649 =  ( n1273____DOLLAR__3173 ) | ( n1462____DOLLAR__3648 )  ;
assign n1464____DOLLAR__3650 =  ( n1272____DOLLAR__3169 ) | ( n1463____DOLLAR__3649 )  ;
assign n1465____DOLLAR__3651 =  ( n1271____DOLLAR__3165 ) | ( n1464____DOLLAR__3650 )  ;
assign n1466____DOLLAR__3652 =  ( n1270____DOLLAR__3161 ) | ( n1465____DOLLAR__3651 )  ;
assign n1467____DOLLAR__3653 =  ( n1269____DOLLAR__3157 ) | ( n1466____DOLLAR__3652 )  ;
assign n1468____DOLLAR__3654 =  ( n1268____DOLLAR__3153 ) | ( n1467____DOLLAR__3653 )  ;
assign n1469____DOLLAR__3655 =  ( n1267____DOLLAR__3149 ) | ( n1468____DOLLAR__3654 )  ;
assign n1470____DOLLAR__3656 =  ( n1266____DOLLAR__3145 ) | ( n1469____DOLLAR__3655 )  ;
assign n1471____DOLLAR__3657 =  ( n1265____DOLLAR__3141 ) | ( n1470____DOLLAR__3656 )  ;
assign n1472____DOLLAR__3658 =  ( n1264____DOLLAR__3137 ) | ( n1471____DOLLAR__3657 )  ;
assign n1473____DOLLAR__3659 =  ( n1263____DOLLAR__3133 ) | ( n1472____DOLLAR__3658 )  ;
assign n1474____DOLLAR__3660 =  ( n1262____DOLLAR__3129 ) | ( n1473____DOLLAR__3659 )  ;
assign n1475____DOLLAR__3661 =  ( n1261____DOLLAR__3125 ) | ( n1474____DOLLAR__3660 )  ;
assign n1476____DOLLAR__3662 =  ( n1260____DOLLAR__3121 ) | ( n1475____DOLLAR__3661 )  ;
assign n1477____DOLLAR__3663 =  ( n1259____DOLLAR__3117 ) | ( n1476____DOLLAR__3662 )  ;
assign n1478____DOLLAR__3664 =  ( n1258____DOLLAR__3113 ) | ( n1477____DOLLAR__3663 )  ;
assign n1479____DOLLAR__3665 =  ( n1257____DOLLAR__3109 ) | ( n1478____DOLLAR__3664 )  ;
assign n1480____DOLLAR__3666 =  ( n1256____DOLLAR__3105 ) | ( n1479____DOLLAR__3665 )  ;
assign n1481____DOLLAR__3667 =  ( n1255____DOLLAR__3101 ) | ( n1480____DOLLAR__3666 )  ;
assign n1482____DOLLAR__3668 =  ( n1254____DOLLAR__3097 ) | ( n1481____DOLLAR__3667 )  ;
assign n1483____DOLLAR__3669 =  ( n1253____DOLLAR__3093 ) | ( n1482____DOLLAR__3668 )  ;
assign n1484____DOLLAR__3670 =  ( n1252____DOLLAR__3089 ) | ( n1483____DOLLAR__3669 )  ;
assign n1485____DOLLAR__3671 =  ( n1251____DOLLAR__3085 ) | ( n1484____DOLLAR__3670 )  ;
assign n1486____DOLLAR__3672 =  ( n1250____DOLLAR__3081 ) | ( n1485____DOLLAR__3671 )  ;
assign n1487____DOLLAR__3673 =  ( n1249____DOLLAR__3077 ) | ( n1486____DOLLAR__3672 )  ;
assign n1488____DOLLAR__3674 =  ( n1248____DOLLAR__3073 ) | ( n1487____DOLLAR__3673 )  ;
assign n1489____DOLLAR__3675 =  ( n1247____DOLLAR__3069 ) | ( n1488____DOLLAR__3674 )  ;
assign n1490____DOLLAR__3676 =  ( n1246____DOLLAR__3065 ) | ( n1489____DOLLAR__3675 )  ;
assign n1491____DOLLAR__3677 =  ( n1245____DOLLAR__3061 ) | ( n1490____DOLLAR__3676 )  ;
assign n1492____DOLLAR__3678 =  ( n1244____DOLLAR__3057 ) | ( n1491____DOLLAR__3677 )  ;
assign n1493____DOLLAR__3679 =  ( n1243____DOLLAR__3053 ) | ( n1492____DOLLAR__3678 )  ;
assign n1494____DOLLAR__3680 =  ( n1242____DOLLAR__3049 ) | ( n1493____DOLLAR__3679 )  ;
assign n1495____DOLLAR__3681 =  ( n1241____DOLLAR__3045 ) | ( n1494____DOLLAR__3680 )  ;
assign n1496____DOLLAR__3682 =  ( n1240____DOLLAR__3041 ) | ( n1495____DOLLAR__3681 )  ;
assign n1497____DOLLAR__3683 =  ( n1239____DOLLAR__3037 ) | ( n1496____DOLLAR__3682 )  ;
assign n1498____DOLLAR__3684 =  ( n1238____DOLLAR__3033 ) | ( n1497____DOLLAR__3683 )  ;
assign n1499____DOLLAR__3685 =  ( n1237____DOLLAR__3029 ) | ( n1498____DOLLAR__3684 )  ;
assign n1500____DOLLAR__3686 =  ( n1236____DOLLAR__3025 ) | ( n1499____DOLLAR__3685 )  ;
assign n1501____DOLLAR__3687 =  ( n1235____DOLLAR__3021 ) | ( n1500____DOLLAR__3686 )  ;
assign n1502____DOLLAR__3688 =  ( n1234____DOLLAR__3017 ) | ( n1501____DOLLAR__3687 )  ;
assign n1503____DOLLAR__3689 =  ( n1233____DOLLAR__3013 ) | ( n1502____DOLLAR__3688 )  ;
assign n1504____DOLLAR__3690 =  ( n1232____DOLLAR__3009 ) | ( n1503____DOLLAR__3689 )  ;
assign n1505____DOLLAR__3691 =  ( n1231____DOLLAR__3005 ) | ( n1504____DOLLAR__3690 )  ;
assign n1506____DOLLAR__3694 =  ( PC ) + ( 16'd1 )  ;
assign n1507____DOLLAR__3695 =  ( n1505____DOLLAR__3691 ) ? ( n1506____DOLLAR__3694 ) : ( PC ) ;
assign n1508____DOLLAR__3696 =  ( n1226____DOLLAR__2976 ) ? ( n1230____DOLLAR__2999 ) : ( n1507____DOLLAR__3695 ) ;
assign n1509____DOLLAR__3697 =  ( n1222____DOLLAR__2949 ) ? ( n1223____DOLLAR__2964 ) : ( n1508____DOLLAR__3696 ) ;
assign n1510____DOLLAR__3698 =  ( n1218____DOLLAR__2935 ) ? ( n1219____DOLLAR__2938 ) : ( n1509____DOLLAR__3697 ) ;
assign n1511____DOLLAR__3699 =  ( n1003____DOLLAR__2462 ) ? ( n1095____DOLLAR__2624 ) : ( n1510____DOLLAR__3698 ) ;
assign n1512____DOLLAR__3700 =  ( n996____DOLLAR__2427 ) ? ( n1000____DOLLAR__2450 ) : ( n1511____DOLLAR__3699 ) ;
assign n1513____DOLLAR__3701 =  ( n925____DOLLAR__2403 ) ? ( n993____DOLLAR__2415 ) : ( n1512____DOLLAR__3700 ) ;
assign n1514____DOLLAR__3706 =  ( oc8051_ROM_rdata_0 ) == ( 8'd255 )  ;
assign n1515____DOLLAR__3710 =  ( oc8051_ROM_rdata_0 ) == ( 8'd254 )  ;
assign n1516____DOLLAR__3714 =  ( oc8051_ROM_rdata_0 ) == ( 8'd253 )  ;
assign n1517____DOLLAR__3718 =  ( oc8051_ROM_rdata_0 ) == ( 8'd252 )  ;
assign n1518____DOLLAR__3722 =  ( oc8051_ROM_rdata_0 ) == ( 8'd251 )  ;
assign n1519____DOLLAR__3726 =  ( oc8051_ROM_rdata_0 ) == ( 8'd250 )  ;
assign n1520____DOLLAR__3730 =  ( oc8051_ROM_rdata_0 ) == ( 8'd249 )  ;
assign n1521____DOLLAR__3734 =  ( oc8051_ROM_rdata_0 ) == ( 8'd248 )  ;
assign n1522____DOLLAR__3738 =  ( oc8051_ROM_rdata_0 ) == ( 8'd247 )  ;
assign n1523____DOLLAR__3742 =  ( oc8051_ROM_rdata_0 ) == ( 8'd246 )  ;
assign n1524____DOLLAR__3746 =  ( oc8051_ROM_rdata_0 ) == ( 8'd244 )  ;
assign n1525____DOLLAR__3750 =  ( oc8051_ROM_rdata_0 ) == ( 8'd243 )  ;
assign n1526____DOLLAR__3754 =  ( oc8051_ROM_rdata_0 ) == ( 8'd242 )  ;
assign n1527____DOLLAR__3758 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign n1528____DOLLAR__3762 =  ( oc8051_ROM_rdata_0 ) == ( 8'd239 )  ;
assign n1529____DOLLAR__3766 =  ( oc8051_ROM_rdata_0 ) == ( 8'd238 )  ;
assign n1530____DOLLAR__3770 =  ( oc8051_ROM_rdata_0 ) == ( 8'd237 )  ;
assign n1531____DOLLAR__3774 =  ( oc8051_ROM_rdata_0 ) == ( 8'd236 )  ;
assign n1532____DOLLAR__3778 =  ( oc8051_ROM_rdata_0 ) == ( 8'd235 )  ;
assign n1533____DOLLAR__3782 =  ( oc8051_ROM_rdata_0 ) == ( 8'd234 )  ;
assign n1534____DOLLAR__3786 =  ( oc8051_ROM_rdata_0 ) == ( 8'd233 )  ;
assign n1535____DOLLAR__3790 =  ( oc8051_ROM_rdata_0 ) == ( 8'd232 )  ;
assign n1536____DOLLAR__3794 =  ( oc8051_ROM_rdata_0 ) == ( 8'd231 )  ;
assign n1537____DOLLAR__3798 =  ( oc8051_ROM_rdata_0 ) == ( 8'd230 )  ;
assign n1538____DOLLAR__3802 =  ( oc8051_ROM_rdata_0 ) == ( 8'd229 )  ;
assign n1539____DOLLAR__3806 =  ( oc8051_ROM_rdata_0 ) == ( 8'd228 )  ;
assign n1540____DOLLAR__3810 =  ( oc8051_ROM_rdata_0 ) == ( 8'd227 )  ;
assign n1541____DOLLAR__3814 =  ( oc8051_ROM_rdata_0 ) == ( 8'd226 )  ;
assign n1542____DOLLAR__3818 =  ( oc8051_ROM_rdata_0 ) == ( 8'd225 )  ;
assign n1543____DOLLAR__3822 =  ( oc8051_ROM_rdata_0 ) == ( 8'd224 )  ;
assign n1544____DOLLAR__3826 =  ( oc8051_ROM_rdata_0 ) == ( 8'd223 )  ;
assign n1545____DOLLAR__3830 =  ( oc8051_ROM_rdata_0 ) == ( 8'd222 )  ;
assign n1546____DOLLAR__3834 =  ( oc8051_ROM_rdata_0 ) == ( 8'd221 )  ;
assign n1547____DOLLAR__3838 =  ( oc8051_ROM_rdata_0 ) == ( 8'd220 )  ;
assign n1548____DOLLAR__3842 =  ( oc8051_ROM_rdata_0 ) == ( 8'd219 )  ;
assign n1549____DOLLAR__3846 =  ( oc8051_ROM_rdata_0 ) == ( 8'd218 )  ;
assign n1550____DOLLAR__3850 =  ( oc8051_ROM_rdata_0 ) == ( 8'd217 )  ;
assign n1551____DOLLAR__3854 =  ( oc8051_ROM_rdata_0 ) == ( 8'd216 )  ;
assign n1552____DOLLAR__3858 =  ( oc8051_ROM_rdata_0 ) == ( 8'd215 )  ;
assign n1553____DOLLAR__3862 =  ( oc8051_ROM_rdata_0 ) == ( 8'd214 )  ;
assign n1554____DOLLAR__3866 =  ( oc8051_ROM_rdata_0 ) == ( 8'd212 )  ;
assign n1555____DOLLAR__3870 =  ( oc8051_ROM_rdata_0 ) == ( 8'd211 )  ;
assign n1556____DOLLAR__3874 =  ( oc8051_ROM_rdata_0 ) == ( 8'd210 )  ;
assign n1557____DOLLAR__3878 =  ( oc8051_ROM_rdata_0 ) == ( 8'd207 )  ;
assign n1558____DOLLAR__3882 =  ( oc8051_ROM_rdata_0 ) == ( 8'd206 )  ;
assign n1559____DOLLAR__3886 =  ( oc8051_ROM_rdata_0 ) == ( 8'd205 )  ;
assign n1560____DOLLAR__3890 =  ( oc8051_ROM_rdata_0 ) == ( 8'd204 )  ;
assign n1561____DOLLAR__3894 =  ( oc8051_ROM_rdata_0 ) == ( 8'd203 )  ;
assign n1562____DOLLAR__3898 =  ( oc8051_ROM_rdata_0 ) == ( 8'd202 )  ;
assign n1563____DOLLAR__3902 =  ( oc8051_ROM_rdata_0 ) == ( 8'd201 )  ;
assign n1564____DOLLAR__3906 =  ( oc8051_ROM_rdata_0 ) == ( 8'd200 )  ;
assign n1565____DOLLAR__3910 =  ( oc8051_ROM_rdata_0 ) == ( 8'd199 )  ;
assign n1566____DOLLAR__3914 =  ( oc8051_ROM_rdata_0 ) == ( 8'd198 )  ;
assign n1567____DOLLAR__3918 =  ( oc8051_ROM_rdata_0 ) == ( 8'd196 )  ;
assign n1568____DOLLAR__3922 =  ( oc8051_ROM_rdata_0 ) == ( 8'd195 )  ;
assign n1569____DOLLAR__3926 =  ( oc8051_ROM_rdata_0 ) == ( 8'd194 )  ;
assign n1570____DOLLAR__3930 =  ( oc8051_ROM_rdata_0 ) == ( 8'd193 )  ;
assign n1571____DOLLAR__3934 =  ( oc8051_ROM_rdata_0 ) == ( 8'd191 )  ;
assign n1572____DOLLAR__3938 =  ( oc8051_ROM_rdata_0 ) == ( 8'd190 )  ;
assign n1573____DOLLAR__3942 =  ( oc8051_ROM_rdata_0 ) == ( 8'd189 )  ;
assign n1574____DOLLAR__3946 =  ( oc8051_ROM_rdata_0 ) == ( 8'd188 )  ;
assign n1575____DOLLAR__3950 =  ( oc8051_ROM_rdata_0 ) == ( 8'd187 )  ;
assign n1576____DOLLAR__3954 =  ( oc8051_ROM_rdata_0 ) == ( 8'd186 )  ;
assign n1577____DOLLAR__3958 =  ( oc8051_ROM_rdata_0 ) == ( 8'd185 )  ;
assign n1578____DOLLAR__3962 =  ( oc8051_ROM_rdata_0 ) == ( 8'd184 )  ;
assign n1579____DOLLAR__3966 =  ( oc8051_ROM_rdata_0 ) == ( 8'd183 )  ;
assign n1580____DOLLAR__3970 =  ( oc8051_ROM_rdata_0 ) == ( 8'd182 )  ;
assign n1581____DOLLAR__3974 =  ( oc8051_ROM_rdata_0 ) == ( 8'd181 )  ;
assign n1582____DOLLAR__3978 =  ( oc8051_ROM_rdata_0 ) == ( 8'd180 )  ;
assign n1583____DOLLAR__3982 =  ( oc8051_ROM_rdata_0 ) == ( 8'd179 )  ;
assign n1584____DOLLAR__3986 =  ( oc8051_ROM_rdata_0 ) == ( 8'd178 )  ;
assign n1585____DOLLAR__3990 =  ( oc8051_ROM_rdata_0 ) == ( 8'd176 )  ;
assign n1586____DOLLAR__3994 =  ( oc8051_ROM_rdata_0 ) == ( 8'd175 )  ;
assign n1587____DOLLAR__3998 =  ( oc8051_ROM_rdata_0 ) == ( 8'd174 )  ;
assign n1588____DOLLAR__4002 =  ( oc8051_ROM_rdata_0 ) == ( 8'd173 )  ;
assign n1589____DOLLAR__4006 =  ( oc8051_ROM_rdata_0 ) == ( 8'd172 )  ;
assign n1590____DOLLAR__4010 =  ( oc8051_ROM_rdata_0 ) == ( 8'd171 )  ;
assign n1591____DOLLAR__4014 =  ( oc8051_ROM_rdata_0 ) == ( 8'd170 )  ;
assign n1592____DOLLAR__4018 =  ( oc8051_ROM_rdata_0 ) == ( 8'd169 )  ;
assign n1593____DOLLAR__4022 =  ( oc8051_ROM_rdata_0 ) == ( 8'd168 )  ;
assign n1594____DOLLAR__4026 =  ( oc8051_ROM_rdata_0 ) == ( 8'd167 )  ;
assign n1595____DOLLAR__4030 =  ( oc8051_ROM_rdata_0 ) == ( 8'd166 )  ;
assign n1596____DOLLAR__4034 =  ( oc8051_ROM_rdata_0 ) == ( 8'd165 )  ;
assign n1597____DOLLAR__4038 =  ( oc8051_ROM_rdata_0 ) == ( 8'd164 )  ;
assign n1598____DOLLAR__4042 =  ( oc8051_ROM_rdata_0 ) == ( 8'd163 )  ;
assign n1599____DOLLAR__4046 =  ( oc8051_ROM_rdata_0 ) == ( 8'd162 )  ;
assign n1600____DOLLAR__4050 =  ( oc8051_ROM_rdata_0 ) == ( 8'd161 )  ;
assign n1601____DOLLAR__4054 =  ( oc8051_ROM_rdata_0 ) == ( 8'd160 )  ;
assign n1602____DOLLAR__4058 =  ( oc8051_ROM_rdata_0 ) == ( 8'd159 )  ;
assign n1603____DOLLAR__4062 =  ( oc8051_ROM_rdata_0 ) == ( 8'd158 )  ;
assign n1604____DOLLAR__4066 =  ( oc8051_ROM_rdata_0 ) == ( 8'd157 )  ;
assign n1605____DOLLAR__4070 =  ( oc8051_ROM_rdata_0 ) == ( 8'd156 )  ;
assign n1606____DOLLAR__4074 =  ( oc8051_ROM_rdata_0 ) == ( 8'd155 )  ;
assign n1607____DOLLAR__4078 =  ( oc8051_ROM_rdata_0 ) == ( 8'd154 )  ;
assign n1608____DOLLAR__4082 =  ( oc8051_ROM_rdata_0 ) == ( 8'd153 )  ;
assign n1609____DOLLAR__4086 =  ( oc8051_ROM_rdata_0 ) == ( 8'd152 )  ;
assign n1610____DOLLAR__4090 =  ( oc8051_ROM_rdata_0 ) == ( 8'd151 )  ;
assign n1611____DOLLAR__4094 =  ( oc8051_ROM_rdata_0 ) == ( 8'd150 )  ;
assign n1612____DOLLAR__4098 =  ( oc8051_ROM_rdata_0 ) == ( 8'd149 )  ;
assign n1613____DOLLAR__4102 =  ( oc8051_ROM_rdata_0 ) == ( 8'd148 )  ;
assign n1614____DOLLAR__4106 =  ( oc8051_ROM_rdata_0 ) == ( 8'd147 )  ;
assign n1615____DOLLAR__4110 =  ( oc8051_ROM_rdata_0 ) == ( 8'd146 )  ;
assign n1616____DOLLAR__4114 =  ( oc8051_ROM_rdata_0 ) == ( 8'd144 )  ;
assign n1617____DOLLAR__4118 =  ( oc8051_ROM_rdata_0 ) == ( 8'd132 )  ;
assign n1618____DOLLAR__4122 =  ( oc8051_ROM_rdata_0 ) == ( 8'd131 )  ;
assign n1619____DOLLAR__4126 =  ( oc8051_ROM_rdata_0 ) == ( 8'd130 )  ;
assign n1620____DOLLAR__4130 =  ( oc8051_ROM_rdata_0 ) == ( 8'd129 )  ;
assign n1621____DOLLAR__4134 =  ( oc8051_ROM_rdata_0 ) == ( 8'd128 )  ;
assign n1622____DOLLAR__4138 =  ( oc8051_ROM_rdata_0 ) == ( 8'd127 )  ;
assign n1623____DOLLAR__4142 =  ( oc8051_ROM_rdata_0 ) == ( 8'd126 )  ;
assign n1624____DOLLAR__4146 =  ( oc8051_ROM_rdata_0 ) == ( 8'd125 )  ;
assign n1625____DOLLAR__4150 =  ( oc8051_ROM_rdata_0 ) == ( 8'd124 )  ;
assign n1626____DOLLAR__4154 =  ( oc8051_ROM_rdata_0 ) == ( 8'd123 )  ;
assign n1627____DOLLAR__4158 =  ( oc8051_ROM_rdata_0 ) == ( 8'd122 )  ;
assign n1628____DOLLAR__4162 =  ( oc8051_ROM_rdata_0 ) == ( 8'd121 )  ;
assign n1629____DOLLAR__4166 =  ( oc8051_ROM_rdata_0 ) == ( 8'd120 )  ;
assign n1630____DOLLAR__4170 =  ( oc8051_ROM_rdata_0 ) == ( 8'd119 )  ;
assign n1631____DOLLAR__4174 =  ( oc8051_ROM_rdata_0 ) == ( 8'd118 )  ;
assign n1632____DOLLAR__4178 =  ( oc8051_ROM_rdata_0 ) == ( 8'd116 )  ;
assign n1633____DOLLAR__4182 =  ( oc8051_ROM_rdata_0 ) == ( 8'd115 )  ;
assign n1634____DOLLAR__4186 =  ( oc8051_ROM_rdata_0 ) == ( 8'd114 )  ;
assign n1635____DOLLAR__4190 =  ( oc8051_ROM_rdata_0 ) == ( 8'd112 )  ;
assign n1636____DOLLAR__4194 =  ( oc8051_ROM_rdata_0 ) == ( 8'd111 )  ;
assign n1637____DOLLAR__4198 =  ( oc8051_ROM_rdata_0 ) == ( 8'd110 )  ;
assign n1638____DOLLAR__4202 =  ( oc8051_ROM_rdata_0 ) == ( 8'd109 )  ;
assign n1639____DOLLAR__4206 =  ( oc8051_ROM_rdata_0 ) == ( 8'd108 )  ;
assign n1640____DOLLAR__4210 =  ( oc8051_ROM_rdata_0 ) == ( 8'd107 )  ;
assign n1641____DOLLAR__4214 =  ( oc8051_ROM_rdata_0 ) == ( 8'd106 )  ;
assign n1642____DOLLAR__4218 =  ( oc8051_ROM_rdata_0 ) == ( 8'd105 )  ;
assign n1643____DOLLAR__4222 =  ( oc8051_ROM_rdata_0 ) == ( 8'd104 )  ;
assign n1644____DOLLAR__4226 =  ( oc8051_ROM_rdata_0 ) == ( 8'd103 )  ;
assign n1645____DOLLAR__4230 =  ( oc8051_ROM_rdata_0 ) == ( 8'd102 )  ;
assign n1646____DOLLAR__4234 =  ( oc8051_ROM_rdata_0 ) == ( 8'd101 )  ;
assign n1647____DOLLAR__4238 =  ( oc8051_ROM_rdata_0 ) == ( 8'd100 )  ;
assign n1648____DOLLAR__4242 =  ( oc8051_ROM_rdata_0 ) == ( 8'd97 )  ;
assign n1649____DOLLAR__4246 =  ( oc8051_ROM_rdata_0 ) == ( 8'd96 )  ;
assign n1650____DOLLAR__4250 =  ( oc8051_ROM_rdata_0 ) == ( 8'd95 )  ;
assign n1651____DOLLAR__4254 =  ( oc8051_ROM_rdata_0 ) == ( 8'd94 )  ;
assign n1652____DOLLAR__4258 =  ( oc8051_ROM_rdata_0 ) == ( 8'd93 )  ;
assign n1653____DOLLAR__4262 =  ( oc8051_ROM_rdata_0 ) == ( 8'd92 )  ;
assign n1654____DOLLAR__4266 =  ( oc8051_ROM_rdata_0 ) == ( 8'd91 )  ;
assign n1655____DOLLAR__4270 =  ( oc8051_ROM_rdata_0 ) == ( 8'd90 )  ;
assign n1656____DOLLAR__4274 =  ( oc8051_ROM_rdata_0 ) == ( 8'd89 )  ;
assign n1657____DOLLAR__4278 =  ( oc8051_ROM_rdata_0 ) == ( 8'd88 )  ;
assign n1658____DOLLAR__4282 =  ( oc8051_ROM_rdata_0 ) == ( 8'd87 )  ;
assign n1659____DOLLAR__4286 =  ( oc8051_ROM_rdata_0 ) == ( 8'd86 )  ;
assign n1660____DOLLAR__4290 =  ( oc8051_ROM_rdata_0 ) == ( 8'd85 )  ;
assign n1661____DOLLAR__4294 =  ( oc8051_ROM_rdata_0 ) == ( 8'd84 )  ;
assign n1662____DOLLAR__4298 =  ( oc8051_ROM_rdata_0 ) == ( 8'd80 )  ;
assign n1663____DOLLAR__4302 =  ( oc8051_ROM_rdata_0 ) == ( 8'd79 )  ;
assign n1664____DOLLAR__4306 =  ( oc8051_ROM_rdata_0 ) == ( 8'd78 )  ;
assign n1665____DOLLAR__4310 =  ( oc8051_ROM_rdata_0 ) == ( 8'd77 )  ;
assign n1666____DOLLAR__4314 =  ( oc8051_ROM_rdata_0 ) == ( 8'd76 )  ;
assign n1667____DOLLAR__4318 =  ( oc8051_ROM_rdata_0 ) == ( 8'd75 )  ;
assign n1668____DOLLAR__4322 =  ( oc8051_ROM_rdata_0 ) == ( 8'd74 )  ;
assign n1669____DOLLAR__4326 =  ( oc8051_ROM_rdata_0 ) == ( 8'd73 )  ;
assign n1670____DOLLAR__4330 =  ( oc8051_ROM_rdata_0 ) == ( 8'd72 )  ;
assign n1671____DOLLAR__4334 =  ( oc8051_ROM_rdata_0 ) == ( 8'd71 )  ;
assign n1672____DOLLAR__4338 =  ( oc8051_ROM_rdata_0 ) == ( 8'd70 )  ;
assign n1673____DOLLAR__4342 =  ( oc8051_ROM_rdata_0 ) == ( 8'd69 )  ;
assign n1674____DOLLAR__4346 =  ( oc8051_ROM_rdata_0 ) == ( 8'd68 )  ;
assign n1675____DOLLAR__4350 =  ( oc8051_ROM_rdata_0 ) == ( 8'd65 )  ;
assign n1676____DOLLAR__4354 =  ( oc8051_ROM_rdata_0 ) == ( 8'd64 )  ;
assign n1677____DOLLAR__4358 =  ( oc8051_ROM_rdata_0 ) == ( 8'd63 )  ;
assign n1678____DOLLAR__4362 =  ( oc8051_ROM_rdata_0 ) == ( 8'd62 )  ;
assign n1679____DOLLAR__4366 =  ( oc8051_ROM_rdata_0 ) == ( 8'd61 )  ;
assign n1680____DOLLAR__4370 =  ( oc8051_ROM_rdata_0 ) == ( 8'd60 )  ;
assign n1681____DOLLAR__4374 =  ( oc8051_ROM_rdata_0 ) == ( 8'd59 )  ;
assign n1682____DOLLAR__4378 =  ( oc8051_ROM_rdata_0 ) == ( 8'd58 )  ;
assign n1683____DOLLAR__4382 =  ( oc8051_ROM_rdata_0 ) == ( 8'd57 )  ;
assign n1684____DOLLAR__4386 =  ( oc8051_ROM_rdata_0 ) == ( 8'd56 )  ;
assign n1685____DOLLAR__4390 =  ( oc8051_ROM_rdata_0 ) == ( 8'd55 )  ;
assign n1686____DOLLAR__4394 =  ( oc8051_ROM_rdata_0 ) == ( 8'd54 )  ;
assign n1687____DOLLAR__4398 =  ( oc8051_ROM_rdata_0 ) == ( 8'd53 )  ;
assign n1688____DOLLAR__4402 =  ( oc8051_ROM_rdata_0 ) == ( 8'd52 )  ;
assign n1689____DOLLAR__4406 =  ( oc8051_ROM_rdata_0 ) == ( 8'd51 )  ;
assign n1690____DOLLAR__4410 =  ( oc8051_ROM_rdata_0 ) == ( 8'd48 )  ;
assign n1691____DOLLAR__4414 =  ( oc8051_ROM_rdata_0 ) == ( 8'd47 )  ;
assign n1692____DOLLAR__4418 =  ( oc8051_ROM_rdata_0 ) == ( 8'd46 )  ;
assign n1693____DOLLAR__4422 =  ( oc8051_ROM_rdata_0 ) == ( 8'd45 )  ;
assign n1694____DOLLAR__4426 =  ( oc8051_ROM_rdata_0 ) == ( 8'd44 )  ;
assign n1695____DOLLAR__4430 =  ( oc8051_ROM_rdata_0 ) == ( 8'd43 )  ;
assign n1696____DOLLAR__4434 =  ( oc8051_ROM_rdata_0 ) == ( 8'd42 )  ;
assign n1697____DOLLAR__4438 =  ( oc8051_ROM_rdata_0 ) == ( 8'd41 )  ;
assign n1698____DOLLAR__4442 =  ( oc8051_ROM_rdata_0 ) == ( 8'd40 )  ;
assign n1699____DOLLAR__4446 =  ( oc8051_ROM_rdata_0 ) == ( 8'd39 )  ;
assign n1700____DOLLAR__4450 =  ( oc8051_ROM_rdata_0 ) == ( 8'd38 )  ;
assign n1701____DOLLAR__4454 =  ( oc8051_ROM_rdata_0 ) == ( 8'd37 )  ;
assign n1702____DOLLAR__4458 =  ( oc8051_ROM_rdata_0 ) == ( 8'd36 )  ;
assign n1703____DOLLAR__4462 =  ( oc8051_ROM_rdata_0 ) == ( 8'd35 )  ;
assign n1704____DOLLAR__4466 =  ( oc8051_ROM_rdata_0 ) == ( 8'd33 )  ;
assign n1705____DOLLAR__4470 =  ( oc8051_ROM_rdata_0 ) == ( 8'd32 )  ;
assign n1706____DOLLAR__4474 =  ( oc8051_ROM_rdata_0 ) == ( 8'd31 )  ;
assign n1707____DOLLAR__4478 =  ( oc8051_ROM_rdata_0 ) == ( 8'd30 )  ;
assign n1708____DOLLAR__4482 =  ( oc8051_ROM_rdata_0 ) == ( 8'd29 )  ;
assign n1709____DOLLAR__4486 =  ( oc8051_ROM_rdata_0 ) == ( 8'd28 )  ;
assign n1710____DOLLAR__4490 =  ( oc8051_ROM_rdata_0 ) == ( 8'd27 )  ;
assign n1711____DOLLAR__4494 =  ( oc8051_ROM_rdata_0 ) == ( 8'd26 )  ;
assign n1712____DOLLAR__4498 =  ( oc8051_ROM_rdata_0 ) == ( 8'd25 )  ;
assign n1713____DOLLAR__4502 =  ( oc8051_ROM_rdata_0 ) == ( 8'd24 )  ;
assign n1714____DOLLAR__4506 =  ( oc8051_ROM_rdata_0 ) == ( 8'd23 )  ;
assign n1715____DOLLAR__4510 =  ( oc8051_ROM_rdata_0 ) == ( 8'd22 )  ;
assign n1716____DOLLAR__4514 =  ( oc8051_ROM_rdata_0 ) == ( 8'd20 )  ;
assign n1717____DOLLAR__4518 =  ( oc8051_ROM_rdata_0 ) == ( 8'd19 )  ;
assign n1718____DOLLAR__4522 =  ( oc8051_ROM_rdata_0 ) == ( 8'd16 )  ;
assign n1719____DOLLAR__4526 =  ( oc8051_ROM_rdata_0 ) == ( 8'd15 )  ;
assign n1720____DOLLAR__4530 =  ( oc8051_ROM_rdata_0 ) == ( 8'd14 )  ;
assign n1721____DOLLAR__4534 =  ( oc8051_ROM_rdata_0 ) == ( 8'd13 )  ;
assign n1722____DOLLAR__4538 =  ( oc8051_ROM_rdata_0 ) == ( 8'd12 )  ;
assign n1723____DOLLAR__4542 =  ( oc8051_ROM_rdata_0 ) == ( 8'd11 )  ;
assign n1724____DOLLAR__4546 =  ( oc8051_ROM_rdata_0 ) == ( 8'd10 )  ;
assign n1725____DOLLAR__4550 =  ( oc8051_ROM_rdata_0 ) == ( 8'd9 )  ;
assign n1726____DOLLAR__4554 =  ( oc8051_ROM_rdata_0 ) == ( 8'd8 )  ;
assign n1727____DOLLAR__4558 =  ( oc8051_ROM_rdata_0 ) == ( 8'd7 )  ;
assign n1728____DOLLAR__4562 =  ( oc8051_ROM_rdata_0 ) == ( 8'd6 )  ;
assign n1729____DOLLAR__4566 =  ( oc8051_ROM_rdata_0 ) == ( 8'd4 )  ;
assign n1730____DOLLAR__4570 =  ( oc8051_ROM_rdata_0 ) == ( 8'd3 )  ;
assign n1731____DOLLAR__4574 =  ( oc8051_ROM_rdata_0 ) == ( 8'd2 )  ;
assign n1732____DOLLAR__4578 =  ( oc8051_ROM_rdata_0 ) == ( 8'd1 )  ;
assign n1733____DOLLAR__4582 =  ( oc8051_ROM_rdata_0 ) == ( 8'd0 )  ;
assign n1734____DOLLAR__4584 =  ( n1732____DOLLAR__4578 ) | ( n1733____DOLLAR__4582 )  ;
assign n1735____DOLLAR__4585 =  ( n1731____DOLLAR__4574 ) | ( n1734____DOLLAR__4584 )  ;
assign n1736____DOLLAR__4586 =  ( n1730____DOLLAR__4570 ) | ( n1735____DOLLAR__4585 )  ;
assign n1737____DOLLAR__4587 =  ( n1729____DOLLAR__4566 ) | ( n1736____DOLLAR__4586 )  ;
assign n1738____DOLLAR__4588 =  ( n1728____DOLLAR__4562 ) | ( n1737____DOLLAR__4587 )  ;
assign n1739____DOLLAR__4589 =  ( n1727____DOLLAR__4558 ) | ( n1738____DOLLAR__4588 )  ;
assign n1740____DOLLAR__4590 =  ( n1726____DOLLAR__4554 ) | ( n1739____DOLLAR__4589 )  ;
assign n1741____DOLLAR__4591 =  ( n1725____DOLLAR__4550 ) | ( n1740____DOLLAR__4590 )  ;
assign n1742____DOLLAR__4592 =  ( n1724____DOLLAR__4546 ) | ( n1741____DOLLAR__4591 )  ;
assign n1743____DOLLAR__4593 =  ( n1723____DOLLAR__4542 ) | ( n1742____DOLLAR__4592 )  ;
assign n1744____DOLLAR__4594 =  ( n1722____DOLLAR__4538 ) | ( n1743____DOLLAR__4593 )  ;
assign n1745____DOLLAR__4595 =  ( n1721____DOLLAR__4534 ) | ( n1744____DOLLAR__4594 )  ;
assign n1746____DOLLAR__4596 =  ( n1720____DOLLAR__4530 ) | ( n1745____DOLLAR__4595 )  ;
assign n1747____DOLLAR__4597 =  ( n1719____DOLLAR__4526 ) | ( n1746____DOLLAR__4596 )  ;
assign n1748____DOLLAR__4598 =  ( n1718____DOLLAR__4522 ) | ( n1747____DOLLAR__4597 )  ;
assign n1749____DOLLAR__4599 =  ( n1717____DOLLAR__4518 ) | ( n1748____DOLLAR__4598 )  ;
assign n1750____DOLLAR__4600 =  ( n1716____DOLLAR__4514 ) | ( n1749____DOLLAR__4599 )  ;
assign n1751____DOLLAR__4601 =  ( n1715____DOLLAR__4510 ) | ( n1750____DOLLAR__4600 )  ;
assign n1752____DOLLAR__4602 =  ( n1714____DOLLAR__4506 ) | ( n1751____DOLLAR__4601 )  ;
assign n1753____DOLLAR__4603 =  ( n1713____DOLLAR__4502 ) | ( n1752____DOLLAR__4602 )  ;
assign n1754____DOLLAR__4604 =  ( n1712____DOLLAR__4498 ) | ( n1753____DOLLAR__4603 )  ;
assign n1755____DOLLAR__4605 =  ( n1711____DOLLAR__4494 ) | ( n1754____DOLLAR__4604 )  ;
assign n1756____DOLLAR__4606 =  ( n1710____DOLLAR__4490 ) | ( n1755____DOLLAR__4605 )  ;
assign n1757____DOLLAR__4607 =  ( n1709____DOLLAR__4486 ) | ( n1756____DOLLAR__4606 )  ;
assign n1758____DOLLAR__4608 =  ( n1708____DOLLAR__4482 ) | ( n1757____DOLLAR__4607 )  ;
assign n1759____DOLLAR__4609 =  ( n1707____DOLLAR__4478 ) | ( n1758____DOLLAR__4608 )  ;
assign n1760____DOLLAR__4610 =  ( n1706____DOLLAR__4474 ) | ( n1759____DOLLAR__4609 )  ;
assign n1761____DOLLAR__4611 =  ( n1705____DOLLAR__4470 ) | ( n1760____DOLLAR__4610 )  ;
assign n1762____DOLLAR__4612 =  ( n1704____DOLLAR__4466 ) | ( n1761____DOLLAR__4611 )  ;
assign n1763____DOLLAR__4613 =  ( n1703____DOLLAR__4462 ) | ( n1762____DOLLAR__4612 )  ;
assign n1764____DOLLAR__4614 =  ( n1702____DOLLAR__4458 ) | ( n1763____DOLLAR__4613 )  ;
assign n1765____DOLLAR__4615 =  ( n1701____DOLLAR__4454 ) | ( n1764____DOLLAR__4614 )  ;
assign n1766____DOLLAR__4616 =  ( n1700____DOLLAR__4450 ) | ( n1765____DOLLAR__4615 )  ;
assign n1767____DOLLAR__4617 =  ( n1699____DOLLAR__4446 ) | ( n1766____DOLLAR__4616 )  ;
assign n1768____DOLLAR__4618 =  ( n1698____DOLLAR__4442 ) | ( n1767____DOLLAR__4617 )  ;
assign n1769____DOLLAR__4619 =  ( n1697____DOLLAR__4438 ) | ( n1768____DOLLAR__4618 )  ;
assign n1770____DOLLAR__4620 =  ( n1696____DOLLAR__4434 ) | ( n1769____DOLLAR__4619 )  ;
assign n1771____DOLLAR__4621 =  ( n1695____DOLLAR__4430 ) | ( n1770____DOLLAR__4620 )  ;
assign n1772____DOLLAR__4622 =  ( n1694____DOLLAR__4426 ) | ( n1771____DOLLAR__4621 )  ;
assign n1773____DOLLAR__4623 =  ( n1693____DOLLAR__4422 ) | ( n1772____DOLLAR__4622 )  ;
assign n1774____DOLLAR__4624 =  ( n1692____DOLLAR__4418 ) | ( n1773____DOLLAR__4623 )  ;
assign n1775____DOLLAR__4625 =  ( n1691____DOLLAR__4414 ) | ( n1774____DOLLAR__4624 )  ;
assign n1776____DOLLAR__4626 =  ( n1690____DOLLAR__4410 ) | ( n1775____DOLLAR__4625 )  ;
assign n1777____DOLLAR__4627 =  ( n1689____DOLLAR__4406 ) | ( n1776____DOLLAR__4626 )  ;
assign n1778____DOLLAR__4628 =  ( n1688____DOLLAR__4402 ) | ( n1777____DOLLAR__4627 )  ;
assign n1779____DOLLAR__4629 =  ( n1687____DOLLAR__4398 ) | ( n1778____DOLLAR__4628 )  ;
assign n1780____DOLLAR__4630 =  ( n1686____DOLLAR__4394 ) | ( n1779____DOLLAR__4629 )  ;
assign n1781____DOLLAR__4631 =  ( n1685____DOLLAR__4390 ) | ( n1780____DOLLAR__4630 )  ;
assign n1782____DOLLAR__4632 =  ( n1684____DOLLAR__4386 ) | ( n1781____DOLLAR__4631 )  ;
assign n1783____DOLLAR__4633 =  ( n1683____DOLLAR__4382 ) | ( n1782____DOLLAR__4632 )  ;
assign n1784____DOLLAR__4634 =  ( n1682____DOLLAR__4378 ) | ( n1783____DOLLAR__4633 )  ;
assign n1785____DOLLAR__4635 =  ( n1681____DOLLAR__4374 ) | ( n1784____DOLLAR__4634 )  ;
assign n1786____DOLLAR__4636 =  ( n1680____DOLLAR__4370 ) | ( n1785____DOLLAR__4635 )  ;
assign n1787____DOLLAR__4637 =  ( n1679____DOLLAR__4366 ) | ( n1786____DOLLAR__4636 )  ;
assign n1788____DOLLAR__4638 =  ( n1678____DOLLAR__4362 ) | ( n1787____DOLLAR__4637 )  ;
assign n1789____DOLLAR__4639 =  ( n1677____DOLLAR__4358 ) | ( n1788____DOLLAR__4638 )  ;
assign n1790____DOLLAR__4640 =  ( n1676____DOLLAR__4354 ) | ( n1789____DOLLAR__4639 )  ;
assign n1791____DOLLAR__4641 =  ( n1675____DOLLAR__4350 ) | ( n1790____DOLLAR__4640 )  ;
assign n1792____DOLLAR__4642 =  ( n1674____DOLLAR__4346 ) | ( n1791____DOLLAR__4641 )  ;
assign n1793____DOLLAR__4643 =  ( n1673____DOLLAR__4342 ) | ( n1792____DOLLAR__4642 )  ;
assign n1794____DOLLAR__4644 =  ( n1672____DOLLAR__4338 ) | ( n1793____DOLLAR__4643 )  ;
assign n1795____DOLLAR__4645 =  ( n1671____DOLLAR__4334 ) | ( n1794____DOLLAR__4644 )  ;
assign n1796____DOLLAR__4646 =  ( n1670____DOLLAR__4330 ) | ( n1795____DOLLAR__4645 )  ;
assign n1797____DOLLAR__4647 =  ( n1669____DOLLAR__4326 ) | ( n1796____DOLLAR__4646 )  ;
assign n1798____DOLLAR__4648 =  ( n1668____DOLLAR__4322 ) | ( n1797____DOLLAR__4647 )  ;
assign n1799____DOLLAR__4649 =  ( n1667____DOLLAR__4318 ) | ( n1798____DOLLAR__4648 )  ;
assign n1800____DOLLAR__4650 =  ( n1666____DOLLAR__4314 ) | ( n1799____DOLLAR__4649 )  ;
assign n1801____DOLLAR__4651 =  ( n1665____DOLLAR__4310 ) | ( n1800____DOLLAR__4650 )  ;
assign n1802____DOLLAR__4652 =  ( n1664____DOLLAR__4306 ) | ( n1801____DOLLAR__4651 )  ;
assign n1803____DOLLAR__4653 =  ( n1663____DOLLAR__4302 ) | ( n1802____DOLLAR__4652 )  ;
assign n1804____DOLLAR__4654 =  ( n1662____DOLLAR__4298 ) | ( n1803____DOLLAR__4653 )  ;
assign n1805____DOLLAR__4655 =  ( n1661____DOLLAR__4294 ) | ( n1804____DOLLAR__4654 )  ;
assign n1806____DOLLAR__4656 =  ( n1660____DOLLAR__4290 ) | ( n1805____DOLLAR__4655 )  ;
assign n1807____DOLLAR__4657 =  ( n1659____DOLLAR__4286 ) | ( n1806____DOLLAR__4656 )  ;
assign n1808____DOLLAR__4658 =  ( n1658____DOLLAR__4282 ) | ( n1807____DOLLAR__4657 )  ;
assign n1809____DOLLAR__4659 =  ( n1657____DOLLAR__4278 ) | ( n1808____DOLLAR__4658 )  ;
assign n1810____DOLLAR__4660 =  ( n1656____DOLLAR__4274 ) | ( n1809____DOLLAR__4659 )  ;
assign n1811____DOLLAR__4661 =  ( n1655____DOLLAR__4270 ) | ( n1810____DOLLAR__4660 )  ;
assign n1812____DOLLAR__4662 =  ( n1654____DOLLAR__4266 ) | ( n1811____DOLLAR__4661 )  ;
assign n1813____DOLLAR__4663 =  ( n1653____DOLLAR__4262 ) | ( n1812____DOLLAR__4662 )  ;
assign n1814____DOLLAR__4664 =  ( n1652____DOLLAR__4258 ) | ( n1813____DOLLAR__4663 )  ;
assign n1815____DOLLAR__4665 =  ( n1651____DOLLAR__4254 ) | ( n1814____DOLLAR__4664 )  ;
assign n1816____DOLLAR__4666 =  ( n1650____DOLLAR__4250 ) | ( n1815____DOLLAR__4665 )  ;
assign n1817____DOLLAR__4667 =  ( n1649____DOLLAR__4246 ) | ( n1816____DOLLAR__4666 )  ;
assign n1818____DOLLAR__4668 =  ( n1648____DOLLAR__4242 ) | ( n1817____DOLLAR__4667 )  ;
assign n1819____DOLLAR__4669 =  ( n1647____DOLLAR__4238 ) | ( n1818____DOLLAR__4668 )  ;
assign n1820____DOLLAR__4670 =  ( n1646____DOLLAR__4234 ) | ( n1819____DOLLAR__4669 )  ;
assign n1821____DOLLAR__4671 =  ( n1645____DOLLAR__4230 ) | ( n1820____DOLLAR__4670 )  ;
assign n1822____DOLLAR__4672 =  ( n1644____DOLLAR__4226 ) | ( n1821____DOLLAR__4671 )  ;
assign n1823____DOLLAR__4673 =  ( n1643____DOLLAR__4222 ) | ( n1822____DOLLAR__4672 )  ;
assign n1824____DOLLAR__4674 =  ( n1642____DOLLAR__4218 ) | ( n1823____DOLLAR__4673 )  ;
assign n1825____DOLLAR__4675 =  ( n1641____DOLLAR__4214 ) | ( n1824____DOLLAR__4674 )  ;
assign n1826____DOLLAR__4676 =  ( n1640____DOLLAR__4210 ) | ( n1825____DOLLAR__4675 )  ;
assign n1827____DOLLAR__4677 =  ( n1639____DOLLAR__4206 ) | ( n1826____DOLLAR__4676 )  ;
assign n1828____DOLLAR__4678 =  ( n1638____DOLLAR__4202 ) | ( n1827____DOLLAR__4677 )  ;
assign n1829____DOLLAR__4679 =  ( n1637____DOLLAR__4198 ) | ( n1828____DOLLAR__4678 )  ;
assign n1830____DOLLAR__4680 =  ( n1636____DOLLAR__4194 ) | ( n1829____DOLLAR__4679 )  ;
assign n1831____DOLLAR__4681 =  ( n1635____DOLLAR__4190 ) | ( n1830____DOLLAR__4680 )  ;
assign n1832____DOLLAR__4682 =  ( n1634____DOLLAR__4186 ) | ( n1831____DOLLAR__4681 )  ;
assign n1833____DOLLAR__4683 =  ( n1633____DOLLAR__4182 ) | ( n1832____DOLLAR__4682 )  ;
assign n1834____DOLLAR__4684 =  ( n1632____DOLLAR__4178 ) | ( n1833____DOLLAR__4683 )  ;
assign n1835____DOLLAR__4685 =  ( n1631____DOLLAR__4174 ) | ( n1834____DOLLAR__4684 )  ;
assign n1836____DOLLAR__4686 =  ( n1630____DOLLAR__4170 ) | ( n1835____DOLLAR__4685 )  ;
assign n1837____DOLLAR__4687 =  ( n1629____DOLLAR__4166 ) | ( n1836____DOLLAR__4686 )  ;
assign n1838____DOLLAR__4688 =  ( n1628____DOLLAR__4162 ) | ( n1837____DOLLAR__4687 )  ;
assign n1839____DOLLAR__4689 =  ( n1627____DOLLAR__4158 ) | ( n1838____DOLLAR__4688 )  ;
assign n1840____DOLLAR__4690 =  ( n1626____DOLLAR__4154 ) | ( n1839____DOLLAR__4689 )  ;
assign n1841____DOLLAR__4691 =  ( n1625____DOLLAR__4150 ) | ( n1840____DOLLAR__4690 )  ;
assign n1842____DOLLAR__4692 =  ( n1624____DOLLAR__4146 ) | ( n1841____DOLLAR__4691 )  ;
assign n1843____DOLLAR__4693 =  ( n1623____DOLLAR__4142 ) | ( n1842____DOLLAR__4692 )  ;
assign n1844____DOLLAR__4694 =  ( n1622____DOLLAR__4138 ) | ( n1843____DOLLAR__4693 )  ;
assign n1845____DOLLAR__4695 =  ( n1621____DOLLAR__4134 ) | ( n1844____DOLLAR__4694 )  ;
assign n1846____DOLLAR__4696 =  ( n1620____DOLLAR__4130 ) | ( n1845____DOLLAR__4695 )  ;
assign n1847____DOLLAR__4697 =  ( n1619____DOLLAR__4126 ) | ( n1846____DOLLAR__4696 )  ;
assign n1848____DOLLAR__4698 =  ( n1618____DOLLAR__4122 ) | ( n1847____DOLLAR__4697 )  ;
assign n1849____DOLLAR__4699 =  ( n1617____DOLLAR__4118 ) | ( n1848____DOLLAR__4698 )  ;
assign n1850____DOLLAR__4700 =  ( n1616____DOLLAR__4114 ) | ( n1849____DOLLAR__4699 )  ;
assign n1851____DOLLAR__4701 =  ( n1615____DOLLAR__4110 ) | ( n1850____DOLLAR__4700 )  ;
assign n1852____DOLLAR__4702 =  ( n1614____DOLLAR__4106 ) | ( n1851____DOLLAR__4701 )  ;
assign n1853____DOLLAR__4703 =  ( n1613____DOLLAR__4102 ) | ( n1852____DOLLAR__4702 )  ;
assign n1854____DOLLAR__4704 =  ( n1612____DOLLAR__4098 ) | ( n1853____DOLLAR__4703 )  ;
assign n1855____DOLLAR__4705 =  ( n1611____DOLLAR__4094 ) | ( n1854____DOLLAR__4704 )  ;
assign n1856____DOLLAR__4706 =  ( n1610____DOLLAR__4090 ) | ( n1855____DOLLAR__4705 )  ;
assign n1857____DOLLAR__4707 =  ( n1609____DOLLAR__4086 ) | ( n1856____DOLLAR__4706 )  ;
assign n1858____DOLLAR__4708 =  ( n1608____DOLLAR__4082 ) | ( n1857____DOLLAR__4707 )  ;
assign n1859____DOLLAR__4709 =  ( n1607____DOLLAR__4078 ) | ( n1858____DOLLAR__4708 )  ;
assign n1860____DOLLAR__4710 =  ( n1606____DOLLAR__4074 ) | ( n1859____DOLLAR__4709 )  ;
assign n1861____DOLLAR__4711 =  ( n1605____DOLLAR__4070 ) | ( n1860____DOLLAR__4710 )  ;
assign n1862____DOLLAR__4712 =  ( n1604____DOLLAR__4066 ) | ( n1861____DOLLAR__4711 )  ;
assign n1863____DOLLAR__4713 =  ( n1603____DOLLAR__4062 ) | ( n1862____DOLLAR__4712 )  ;
assign n1864____DOLLAR__4714 =  ( n1602____DOLLAR__4058 ) | ( n1863____DOLLAR__4713 )  ;
assign n1865____DOLLAR__4715 =  ( n1601____DOLLAR__4054 ) | ( n1864____DOLLAR__4714 )  ;
assign n1866____DOLLAR__4716 =  ( n1600____DOLLAR__4050 ) | ( n1865____DOLLAR__4715 )  ;
assign n1867____DOLLAR__4717 =  ( n1599____DOLLAR__4046 ) | ( n1866____DOLLAR__4716 )  ;
assign n1868____DOLLAR__4718 =  ( n1598____DOLLAR__4042 ) | ( n1867____DOLLAR__4717 )  ;
assign n1869____DOLLAR__4719 =  ( n1597____DOLLAR__4038 ) | ( n1868____DOLLAR__4718 )  ;
assign n1870____DOLLAR__4720 =  ( n1596____DOLLAR__4034 ) | ( n1869____DOLLAR__4719 )  ;
assign n1871____DOLLAR__4721 =  ( n1595____DOLLAR__4030 ) | ( n1870____DOLLAR__4720 )  ;
assign n1872____DOLLAR__4722 =  ( n1594____DOLLAR__4026 ) | ( n1871____DOLLAR__4721 )  ;
assign n1873____DOLLAR__4723 =  ( n1593____DOLLAR__4022 ) | ( n1872____DOLLAR__4722 )  ;
assign n1874____DOLLAR__4724 =  ( n1592____DOLLAR__4018 ) | ( n1873____DOLLAR__4723 )  ;
assign n1875____DOLLAR__4725 =  ( n1591____DOLLAR__4014 ) | ( n1874____DOLLAR__4724 )  ;
assign n1876____DOLLAR__4726 =  ( n1590____DOLLAR__4010 ) | ( n1875____DOLLAR__4725 )  ;
assign n1877____DOLLAR__4727 =  ( n1589____DOLLAR__4006 ) | ( n1876____DOLLAR__4726 )  ;
assign n1878____DOLLAR__4728 =  ( n1588____DOLLAR__4002 ) | ( n1877____DOLLAR__4727 )  ;
assign n1879____DOLLAR__4729 =  ( n1587____DOLLAR__3998 ) | ( n1878____DOLLAR__4728 )  ;
assign n1880____DOLLAR__4730 =  ( n1586____DOLLAR__3994 ) | ( n1879____DOLLAR__4729 )  ;
assign n1881____DOLLAR__4731 =  ( n1585____DOLLAR__3990 ) | ( n1880____DOLLAR__4730 )  ;
assign n1882____DOLLAR__4732 =  ( n1584____DOLLAR__3986 ) | ( n1881____DOLLAR__4731 )  ;
assign n1883____DOLLAR__4733 =  ( n1583____DOLLAR__3982 ) | ( n1882____DOLLAR__4732 )  ;
assign n1884____DOLLAR__4734 =  ( n1582____DOLLAR__3978 ) | ( n1883____DOLLAR__4733 )  ;
assign n1885____DOLLAR__4735 =  ( n1581____DOLLAR__3974 ) | ( n1884____DOLLAR__4734 )  ;
assign n1886____DOLLAR__4736 =  ( n1580____DOLLAR__3970 ) | ( n1885____DOLLAR__4735 )  ;
assign n1887____DOLLAR__4737 =  ( n1579____DOLLAR__3966 ) | ( n1886____DOLLAR__4736 )  ;
assign n1888____DOLLAR__4738 =  ( n1578____DOLLAR__3962 ) | ( n1887____DOLLAR__4737 )  ;
assign n1889____DOLLAR__4739 =  ( n1577____DOLLAR__3958 ) | ( n1888____DOLLAR__4738 )  ;
assign n1890____DOLLAR__4740 =  ( n1576____DOLLAR__3954 ) | ( n1889____DOLLAR__4739 )  ;
assign n1891____DOLLAR__4741 =  ( n1575____DOLLAR__3950 ) | ( n1890____DOLLAR__4740 )  ;
assign n1892____DOLLAR__4742 =  ( n1574____DOLLAR__3946 ) | ( n1891____DOLLAR__4741 )  ;
assign n1893____DOLLAR__4743 =  ( n1573____DOLLAR__3942 ) | ( n1892____DOLLAR__4742 )  ;
assign n1894____DOLLAR__4744 =  ( n1572____DOLLAR__3938 ) | ( n1893____DOLLAR__4743 )  ;
assign n1895____DOLLAR__4745 =  ( n1571____DOLLAR__3934 ) | ( n1894____DOLLAR__4744 )  ;
assign n1896____DOLLAR__4746 =  ( n1570____DOLLAR__3930 ) | ( n1895____DOLLAR__4745 )  ;
assign n1897____DOLLAR__4747 =  ( n1569____DOLLAR__3926 ) | ( n1896____DOLLAR__4746 )  ;
assign n1898____DOLLAR__4748 =  ( n1568____DOLLAR__3922 ) | ( n1897____DOLLAR__4747 )  ;
assign n1899____DOLLAR__4749 =  ( n1567____DOLLAR__3918 ) | ( n1898____DOLLAR__4748 )  ;
assign n1900____DOLLAR__4750 =  ( n1566____DOLLAR__3914 ) | ( n1899____DOLLAR__4749 )  ;
assign n1901____DOLLAR__4751 =  ( n1565____DOLLAR__3910 ) | ( n1900____DOLLAR__4750 )  ;
assign n1902____DOLLAR__4752 =  ( n1564____DOLLAR__3906 ) | ( n1901____DOLLAR__4751 )  ;
assign n1903____DOLLAR__4753 =  ( n1563____DOLLAR__3902 ) | ( n1902____DOLLAR__4752 )  ;
assign n1904____DOLLAR__4754 =  ( n1562____DOLLAR__3898 ) | ( n1903____DOLLAR__4753 )  ;
assign n1905____DOLLAR__4755 =  ( n1561____DOLLAR__3894 ) | ( n1904____DOLLAR__4754 )  ;
assign n1906____DOLLAR__4756 =  ( n1560____DOLLAR__3890 ) | ( n1905____DOLLAR__4755 )  ;
assign n1907____DOLLAR__4757 =  ( n1559____DOLLAR__3886 ) | ( n1906____DOLLAR__4756 )  ;
assign n1908____DOLLAR__4758 =  ( n1558____DOLLAR__3882 ) | ( n1907____DOLLAR__4757 )  ;
assign n1909____DOLLAR__4759 =  ( n1557____DOLLAR__3878 ) | ( n1908____DOLLAR__4758 )  ;
assign n1910____DOLLAR__4760 =  ( n1556____DOLLAR__3874 ) | ( n1909____DOLLAR__4759 )  ;
assign n1911____DOLLAR__4761 =  ( n1555____DOLLAR__3870 ) | ( n1910____DOLLAR__4760 )  ;
assign n1912____DOLLAR__4762 =  ( n1554____DOLLAR__3866 ) | ( n1911____DOLLAR__4761 )  ;
assign n1913____DOLLAR__4763 =  ( n1553____DOLLAR__3862 ) | ( n1912____DOLLAR__4762 )  ;
assign n1914____DOLLAR__4764 =  ( n1552____DOLLAR__3858 ) | ( n1913____DOLLAR__4763 )  ;
assign n1915____DOLLAR__4765 =  ( n1551____DOLLAR__3854 ) | ( n1914____DOLLAR__4764 )  ;
assign n1916____DOLLAR__4766 =  ( n1550____DOLLAR__3850 ) | ( n1915____DOLLAR__4765 )  ;
assign n1917____DOLLAR__4767 =  ( n1549____DOLLAR__3846 ) | ( n1916____DOLLAR__4766 )  ;
assign n1918____DOLLAR__4768 =  ( n1548____DOLLAR__3842 ) | ( n1917____DOLLAR__4767 )  ;
assign n1919____DOLLAR__4769 =  ( n1547____DOLLAR__3838 ) | ( n1918____DOLLAR__4768 )  ;
assign n1920____DOLLAR__4770 =  ( n1546____DOLLAR__3834 ) | ( n1919____DOLLAR__4769 )  ;
assign n1921____DOLLAR__4771 =  ( n1545____DOLLAR__3830 ) | ( n1920____DOLLAR__4770 )  ;
assign n1922____DOLLAR__4772 =  ( n1544____DOLLAR__3826 ) | ( n1921____DOLLAR__4771 )  ;
assign n1923____DOLLAR__4773 =  ( n1543____DOLLAR__3822 ) | ( n1922____DOLLAR__4772 )  ;
assign n1924____DOLLAR__4774 =  ( n1542____DOLLAR__3818 ) | ( n1923____DOLLAR__4773 )  ;
assign n1925____DOLLAR__4775 =  ( n1541____DOLLAR__3814 ) | ( n1924____DOLLAR__4774 )  ;
assign n1926____DOLLAR__4776 =  ( n1540____DOLLAR__3810 ) | ( n1925____DOLLAR__4775 )  ;
assign n1927____DOLLAR__4777 =  ( n1539____DOLLAR__3806 ) | ( n1926____DOLLAR__4776 )  ;
assign n1928____DOLLAR__4778 =  ( n1538____DOLLAR__3802 ) | ( n1927____DOLLAR__4777 )  ;
assign n1929____DOLLAR__4779 =  ( n1537____DOLLAR__3798 ) | ( n1928____DOLLAR__4778 )  ;
assign n1930____DOLLAR__4780 =  ( n1536____DOLLAR__3794 ) | ( n1929____DOLLAR__4779 )  ;
assign n1931____DOLLAR__4781 =  ( n1535____DOLLAR__3790 ) | ( n1930____DOLLAR__4780 )  ;
assign n1932____DOLLAR__4782 =  ( n1534____DOLLAR__3786 ) | ( n1931____DOLLAR__4781 )  ;
assign n1933____DOLLAR__4783 =  ( n1533____DOLLAR__3782 ) | ( n1932____DOLLAR__4782 )  ;
assign n1934____DOLLAR__4784 =  ( n1532____DOLLAR__3778 ) | ( n1933____DOLLAR__4783 )  ;
assign n1935____DOLLAR__4785 =  ( n1531____DOLLAR__3774 ) | ( n1934____DOLLAR__4784 )  ;
assign n1936____DOLLAR__4786 =  ( n1530____DOLLAR__3770 ) | ( n1935____DOLLAR__4785 )  ;
assign n1937____DOLLAR__4787 =  ( n1529____DOLLAR__3766 ) | ( n1936____DOLLAR__4786 )  ;
assign n1938____DOLLAR__4788 =  ( n1528____DOLLAR__3762 ) | ( n1937____DOLLAR__4787 )  ;
assign n1939____DOLLAR__4789 =  ( n1527____DOLLAR__3758 ) | ( n1938____DOLLAR__4788 )  ;
assign n1940____DOLLAR__4790 =  ( n1526____DOLLAR__3754 ) | ( n1939____DOLLAR__4789 )  ;
assign n1941____DOLLAR__4791 =  ( n1525____DOLLAR__3750 ) | ( n1940____DOLLAR__4790 )  ;
assign n1942____DOLLAR__4792 =  ( n1524____DOLLAR__3746 ) | ( n1941____DOLLAR__4791 )  ;
assign n1943____DOLLAR__4793 =  ( n1523____DOLLAR__3742 ) | ( n1942____DOLLAR__4792 )  ;
assign n1944____DOLLAR__4794 =  ( n1522____DOLLAR__3738 ) | ( n1943____DOLLAR__4793 )  ;
assign n1945____DOLLAR__4795 =  ( n1521____DOLLAR__3734 ) | ( n1944____DOLLAR__4794 )  ;
assign n1946____DOLLAR__4796 =  ( n1520____DOLLAR__3730 ) | ( n1945____DOLLAR__4795 )  ;
assign n1947____DOLLAR__4797 =  ( n1519____DOLLAR__3726 ) | ( n1946____DOLLAR__4796 )  ;
assign n1948____DOLLAR__4798 =  ( n1518____DOLLAR__3722 ) | ( n1947____DOLLAR__4797 )  ;
assign n1949____DOLLAR__4799 =  ( n1517____DOLLAR__3718 ) | ( n1948____DOLLAR__4798 )  ;
assign n1950____DOLLAR__4800 =  ( n1516____DOLLAR__3714 ) | ( n1949____DOLLAR__4799 )  ;
assign n1951____DOLLAR__4801 =  ( n1515____DOLLAR__3710 ) | ( n1950____DOLLAR__4800 )  ;
assign n1952____DOLLAR__4802 =  ( n1514____DOLLAR__3706 ) | ( n1951____DOLLAR__4801 )  ;
assign n1953____DOLLAR__4808 = oc8051_ROM_rdata_1[7:7] ;
assign n1954____DOLLAR__4812 =  ( n1953____DOLLAR__4808 ) == ( 1'd1 )  ;
assign n1955____DOLLAR__4814 = oc8051_ROM_rdata_1[7:3] ;
assign n1956____DOLLAR__4822 =  { ( n1955____DOLLAR__4814 ) , ( 3'd0 ) }  ;
assign n1957____DOLLAR__4824 =  {3'd0 , n1955____DOLLAR__4814}  ;
assign n1958____DOLLAR__4828 =  ( n1957____DOLLAR__4824 ) + ( 8'd32 )  ;
assign n1959____DOLLAR__4829 =  ( n1954____DOLLAR__4812 ) ? ( n1956____DOLLAR__4822 ) : ( n1958____DOLLAR__4828 ) ;
assign n1960____DOLLAR__4832 =  ( n1959____DOLLAR__4829 ) == ( 8'd129 )  ;
assign n1961____DOLLAR__4839 = oc8051_ROM_rdata_1[2:0] ;
assign n1962____DOLLAR__4841 =  {5'd0 , n1961____DOLLAR__4839}  ;
assign n1963____DOLLAR__4843 =  ( 8'd1 ) << ( n1962____DOLLAR__4841 )  ;
assign n1964____DOLLAR__4844 = ~ ( n1963____DOLLAR__4843 ) ;
assign n1965____DOLLAR__4848 = oc8051_ROM_rdata_1[7:7] ;
assign n1966____DOLLAR__4850 =  ( n1965____DOLLAR__4848 ) == ( 1'd1 )  ;
assign n1967____DOLLAR__4852 = oc8051_ROM_rdata_1[7:3] ;
assign n1968____DOLLAR__4858 =  { ( n1967____DOLLAR__4852 ) , ( 3'd0 ) }  ;
assign n1969____DOLLAR__4860 =  {3'd0 , n1967____DOLLAR__4852}  ;
assign n1970____DOLLAR__4862 =  ( n1969____DOLLAR__4860 ) + ( 8'd32 )  ;
assign n1971____DOLLAR__4863 =  ( n1966____DOLLAR__4850 ) ? ( n1968____DOLLAR__4858 ) : ( n1970____DOLLAR__4862 ) ;
assign n1972____DOLLAR__4864 = n1971____DOLLAR__4863[7:7] ;
assign n1973____DOLLAR__4868 =  ( n1972____DOLLAR__4864 ) == ( 1'd0 )  ;
assign n1974____DOLLAR__4873 = oc8051_ROM_rdata_1[7:7] ;
assign n1975____DOLLAR__4875 =  ( n1974____DOLLAR__4873 ) == ( 1'd1 )  ;
assign n1976____DOLLAR__4880 = oc8051_ROM_rdata_1[7:3] ;
assign n1977____DOLLAR__4886 =  { ( n1976____DOLLAR__4880 ) , ( 3'd0 ) }  ;
assign n1978____DOLLAR__4891 = oc8051_ROM_rdata_1[7:3] ;
assign n1979____DOLLAR__4893 =  {3'd0 , n1978____DOLLAR__4891}  ;
assign n1980____DOLLAR__4895 =  ( n1979____DOLLAR__4893 ) + ( 8'd32 )  ;
assign n1981____DOLLAR__4896 =  ( n1975____DOLLAR__4875 ) ? ( n1977____DOLLAR__4886 ) : ( n1980____DOLLAR__4895 ) ;
assign n1982____DOLLAR__187085 = n1981____DOLLAR__4896[3:0] ;
assign n1983____DOLLAR__187166 =  ( n1982____DOLLAR__187085 ) == ( 4'd15 )  ;
assign n1984____DOLLAR__187161 =  ( n1982____DOLLAR__187085 ) == ( 4'd14 )  ;
assign n1985____DOLLAR__187156 =  ( n1982____DOLLAR__187085 ) == ( 4'd13 )  ;
assign n1986____DOLLAR__187151 =  ( n1982____DOLLAR__187085 ) == ( 4'd12 )  ;
assign n1987____DOLLAR__187146 =  ( n1982____DOLLAR__187085 ) == ( 4'd11 )  ;
assign n1988____DOLLAR__187141 =  ( n1982____DOLLAR__187085 ) == ( 4'd10 )  ;
assign n1989____DOLLAR__187136 =  ( n1982____DOLLAR__187085 ) == ( 4'd9 )  ;
assign n1990____DOLLAR__187131 =  ( n1982____DOLLAR__187085 ) == ( 4'd8 )  ;
assign n1991____DOLLAR__187126 =  ( n1982____DOLLAR__187085 ) == ( 4'd7 )  ;
assign n1992____DOLLAR__187121 =  ( n1982____DOLLAR__187085 ) == ( 4'd6 )  ;
assign n1993____DOLLAR__187116 =  ( n1982____DOLLAR__187085 ) == ( 4'd5 )  ;
assign n1994____DOLLAR__187111 =  ( n1982____DOLLAR__187085 ) == ( 4'd4 )  ;
assign n1995____DOLLAR__187106 =  ( n1982____DOLLAR__187085 ) == ( 4'd3 )  ;
assign n1996____DOLLAR__187101 =  ( n1982____DOLLAR__187085 ) == ( 4'd2 )  ;
assign n1997____DOLLAR__187096 =  ( n1982____DOLLAR__187085 ) == ( 4'd1 )  ;
assign n1998____DOLLAR__187091 =  ( n1982____DOLLAR__187085 ) == ( 4'd0 )  ;
assign n1999____DOLLAR__187093 =  ( n1998____DOLLAR__187091 ) ? ( oc8051_IRAM_data_0 ) : ( 8'd0 ) ;
assign n2000____DOLLAR__187098 =  ( n1997____DOLLAR__187096 ) ? ( oc8051_IRAM_data_1 ) : ( n1999____DOLLAR__187093 ) ;
assign n2001____DOLLAR__187103 =  ( n1996____DOLLAR__187101 ) ? ( oc8051_IRAM_data_2 ) : ( n2000____DOLLAR__187098 ) ;
assign n2002____DOLLAR__187108 =  ( n1995____DOLLAR__187106 ) ? ( oc8051_IRAM_data_3 ) : ( n2001____DOLLAR__187103 ) ;
assign n2003____DOLLAR__187113 =  ( n1994____DOLLAR__187111 ) ? ( oc8051_IRAM_data_4 ) : ( n2002____DOLLAR__187108 ) ;
assign n2004____DOLLAR__187118 =  ( n1993____DOLLAR__187116 ) ? ( oc8051_IRAM_data_5 ) : ( n2003____DOLLAR__187113 ) ;
assign n2005____DOLLAR__187123 =  ( n1992____DOLLAR__187121 ) ? ( oc8051_IRAM_data_6 ) : ( n2004____DOLLAR__187118 ) ;
assign n2006____DOLLAR__187128 =  ( n1991____DOLLAR__187126 ) ? ( oc8051_IRAM_data_7 ) : ( n2005____DOLLAR__187123 ) ;
assign n2007____DOLLAR__187133 =  ( n1990____DOLLAR__187131 ) ? ( oc8051_IRAM_data_8 ) : ( n2006____DOLLAR__187128 ) ;
assign n2008____DOLLAR__187138 =  ( n1989____DOLLAR__187136 ) ? ( oc8051_IRAM_data_9 ) : ( n2007____DOLLAR__187133 ) ;
assign n2009____DOLLAR__187143 =  ( n1988____DOLLAR__187141 ) ? ( oc8051_IRAM_data_10 ) : ( n2008____DOLLAR__187138 ) ;
assign n2010____DOLLAR__187148 =  ( n1987____DOLLAR__187146 ) ? ( oc8051_IRAM_data_11 ) : ( n2009____DOLLAR__187143 ) ;
assign n2011____DOLLAR__187153 =  ( n1986____DOLLAR__187151 ) ? ( oc8051_IRAM_data_12 ) : ( n2010____DOLLAR__187148 ) ;
assign n2012____DOLLAR__187158 =  ( n1985____DOLLAR__187156 ) ? ( oc8051_IRAM_data_13 ) : ( n2011____DOLLAR__187153 ) ;
assign n2013____DOLLAR__187163 =  ( n1984____DOLLAR__187161 ) ? ( oc8051_IRAM_data_14 ) : ( n2012____DOLLAR__187158 ) ;
assign n2014____DOLLAR__187168 =  ( n1983____DOLLAR__187166 ) ? ( oc8051_IRAM_data_15 ) : ( n2013____DOLLAR__187163 ) ;
assign n2015____DOLLAR__4902 = oc8051_ROM_rdata_1[7:7] ;
assign n2016____DOLLAR__4904 =  ( n2015____DOLLAR__4902 ) == ( 1'd1 )  ;
assign n2017____DOLLAR__4906 = oc8051_ROM_rdata_1[7:3] ;
assign n2018____DOLLAR__4912 =  { ( n2017____DOLLAR__4906 ) , ( 3'd0 ) }  ;
assign n2019____DOLLAR__4914 =  {3'd0 , n2017____DOLLAR__4906}  ;
assign n2020____DOLLAR__4916 =  ( n2019____DOLLAR__4914 ) + ( 8'd32 )  ;
assign n2021____DOLLAR__4917 =  ( n2016____DOLLAR__4904 ) ? ( n2018____DOLLAR__4912 ) : ( n2020____DOLLAR__4916 ) ;
assign n2022____DOLLAR__4920 =  ( n2021____DOLLAR__4917 ) == ( 8'd128 )  ;
assign n2023____DOLLAR__4925 = oc8051_ROM_rdata_1[7:7] ;
assign n2024____DOLLAR__4927 =  ( n2023____DOLLAR__4925 ) == ( 1'd1 )  ;
assign n2025____DOLLAR__4929 = oc8051_ROM_rdata_1[7:3] ;
assign n2026____DOLLAR__4935 =  { ( n2025____DOLLAR__4929 ) , ( 3'd0 ) }  ;
assign n2027____DOLLAR__4937 =  {3'd0 , n2025____DOLLAR__4929}  ;
assign n2028____DOLLAR__4939 =  ( n2027____DOLLAR__4937 ) + ( 8'd32 )  ;
assign n2029____DOLLAR__4940 =  ( n2024____DOLLAR__4927 ) ? ( n2026____DOLLAR__4935 ) : ( n2028____DOLLAR__4939 ) ;
assign n2030____DOLLAR__4943 =  ( n2029____DOLLAR__4940 ) == ( 8'd129 )  ;
assign n2031____DOLLAR__4948 = oc8051_ROM_rdata_1[7:7] ;
assign n2032____DOLLAR__4950 =  ( n2031____DOLLAR__4948 ) == ( 1'd1 )  ;
assign n2033____DOLLAR__4952 = oc8051_ROM_rdata_1[7:3] ;
assign n2034____DOLLAR__4958 =  { ( n2033____DOLLAR__4952 ) , ( 3'd0 ) }  ;
assign n2035____DOLLAR__4960 =  {3'd0 , n2033____DOLLAR__4952}  ;
assign n2036____DOLLAR__4962 =  ( n2035____DOLLAR__4960 ) + ( 8'd32 )  ;
assign n2037____DOLLAR__4963 =  ( n2032____DOLLAR__4950 ) ? ( n2034____DOLLAR__4958 ) : ( n2036____DOLLAR__4962 ) ;
assign n2038____DOLLAR__4966 =  ( n2037____DOLLAR__4963 ) == ( 8'd130 )  ;
assign n2039____DOLLAR__4971 = oc8051_ROM_rdata_1[7:7] ;
assign n2040____DOLLAR__4973 =  ( n2039____DOLLAR__4971 ) == ( 1'd1 )  ;
assign n2041____DOLLAR__4975 = oc8051_ROM_rdata_1[7:3] ;
assign n2042____DOLLAR__4981 =  { ( n2041____DOLLAR__4975 ) , ( 3'd0 ) }  ;
assign n2043____DOLLAR__4983 =  {3'd0 , n2041____DOLLAR__4975}  ;
assign n2044____DOLLAR__4985 =  ( n2043____DOLLAR__4983 ) + ( 8'd32 )  ;
assign n2045____DOLLAR__4986 =  ( n2040____DOLLAR__4973 ) ? ( n2042____DOLLAR__4981 ) : ( n2044____DOLLAR__4985 ) ;
assign n2046____DOLLAR__4989 =  ( n2045____DOLLAR__4986 ) == ( 8'd131 )  ;
assign n2047____DOLLAR__4994 = oc8051_ROM_rdata_1[7:7] ;
assign n2048____DOLLAR__4996 =  ( n2047____DOLLAR__4994 ) == ( 1'd1 )  ;
assign n2049____DOLLAR__4998 = oc8051_ROM_rdata_1[7:3] ;
assign n2050____DOLLAR__5004 =  { ( n2049____DOLLAR__4998 ) , ( 3'd0 ) }  ;
assign n2051____DOLLAR__5006 =  {3'd0 , n2049____DOLLAR__4998}  ;
assign n2052____DOLLAR__5008 =  ( n2051____DOLLAR__5006 ) + ( 8'd32 )  ;
assign n2053____DOLLAR__5009 =  ( n2048____DOLLAR__4996 ) ? ( n2050____DOLLAR__5004 ) : ( n2052____DOLLAR__5008 ) ;
assign n2054____DOLLAR__5012 =  ( n2053____DOLLAR__5009 ) == ( 8'd135 )  ;
assign n2055____DOLLAR__5017 = oc8051_ROM_rdata_1[7:7] ;
assign n2056____DOLLAR__5019 =  ( n2055____DOLLAR__5017 ) == ( 1'd1 )  ;
assign n2057____DOLLAR__5021 = oc8051_ROM_rdata_1[7:3] ;
assign n2058____DOLLAR__5027 =  { ( n2057____DOLLAR__5021 ) , ( 3'd0 ) }  ;
assign n2059____DOLLAR__5029 =  {3'd0 , n2057____DOLLAR__5021}  ;
assign n2060____DOLLAR__5031 =  ( n2059____DOLLAR__5029 ) + ( 8'd32 )  ;
assign n2061____DOLLAR__5032 =  ( n2056____DOLLAR__5019 ) ? ( n2058____DOLLAR__5027 ) : ( n2060____DOLLAR__5031 ) ;
assign n2062____DOLLAR__5035 =  ( n2061____DOLLAR__5032 ) == ( 8'd136 )  ;
assign n2063____DOLLAR__5040 = oc8051_ROM_rdata_1[7:7] ;
assign n2064____DOLLAR__5042 =  ( n2063____DOLLAR__5040 ) == ( 1'd1 )  ;
assign n2065____DOLLAR__5044 = oc8051_ROM_rdata_1[7:3] ;
assign n2066____DOLLAR__5050 =  { ( n2065____DOLLAR__5044 ) , ( 3'd0 ) }  ;
assign n2067____DOLLAR__5052 =  {3'd0 , n2065____DOLLAR__5044}  ;
assign n2068____DOLLAR__5054 =  ( n2067____DOLLAR__5052 ) + ( 8'd32 )  ;
assign n2069____DOLLAR__5055 =  ( n2064____DOLLAR__5042 ) ? ( n2066____DOLLAR__5050 ) : ( n2068____DOLLAR__5054 ) ;
assign n2070____DOLLAR__5058 =  ( n2069____DOLLAR__5055 ) == ( 8'd137 )  ;
assign n2071____DOLLAR__5063 = oc8051_ROM_rdata_1[7:7] ;
assign n2072____DOLLAR__5065 =  ( n2071____DOLLAR__5063 ) == ( 1'd1 )  ;
assign n2073____DOLLAR__5067 = oc8051_ROM_rdata_1[7:3] ;
assign n2074____DOLLAR__5073 =  { ( n2073____DOLLAR__5067 ) , ( 3'd0 ) }  ;
assign n2075____DOLLAR__5075 =  {3'd0 , n2073____DOLLAR__5067}  ;
assign n2076____DOLLAR__5077 =  ( n2075____DOLLAR__5075 ) + ( 8'd32 )  ;
assign n2077____DOLLAR__5078 =  ( n2072____DOLLAR__5065 ) ? ( n2074____DOLLAR__5073 ) : ( n2076____DOLLAR__5077 ) ;
assign n2078____DOLLAR__5081 =  ( n2077____DOLLAR__5078 ) == ( 8'd138 )  ;
assign n2079____DOLLAR__5086 = oc8051_ROM_rdata_1[7:7] ;
assign n2080____DOLLAR__5088 =  ( n2079____DOLLAR__5086 ) == ( 1'd1 )  ;
assign n2081____DOLLAR__5090 = oc8051_ROM_rdata_1[7:3] ;
assign n2082____DOLLAR__5096 =  { ( n2081____DOLLAR__5090 ) , ( 3'd0 ) }  ;
assign n2083____DOLLAR__5098 =  {3'd0 , n2081____DOLLAR__5090}  ;
assign n2084____DOLLAR__5100 =  ( n2083____DOLLAR__5098 ) + ( 8'd32 )  ;
assign n2085____DOLLAR__5101 =  ( n2080____DOLLAR__5088 ) ? ( n2082____DOLLAR__5096 ) : ( n2084____DOLLAR__5100 ) ;
assign n2086____DOLLAR__5104 =  ( n2085____DOLLAR__5101 ) == ( 8'd140 )  ;
assign n2087____DOLLAR__5109 = oc8051_ROM_rdata_1[7:7] ;
assign n2088____DOLLAR__5111 =  ( n2087____DOLLAR__5109 ) == ( 1'd1 )  ;
assign n2089____DOLLAR__5113 = oc8051_ROM_rdata_1[7:3] ;
assign n2090____DOLLAR__5119 =  { ( n2089____DOLLAR__5113 ) , ( 3'd0 ) }  ;
assign n2091____DOLLAR__5121 =  {3'd0 , n2089____DOLLAR__5113}  ;
assign n2092____DOLLAR__5123 =  ( n2091____DOLLAR__5121 ) + ( 8'd32 )  ;
assign n2093____DOLLAR__5124 =  ( n2088____DOLLAR__5111 ) ? ( n2090____DOLLAR__5119 ) : ( n2092____DOLLAR__5123 ) ;
assign n2094____DOLLAR__5127 =  ( n2093____DOLLAR__5124 ) == ( 8'd139 )  ;
assign n2095____DOLLAR__5132 = oc8051_ROM_rdata_1[7:7] ;
assign n2096____DOLLAR__5134 =  ( n2095____DOLLAR__5132 ) == ( 1'd1 )  ;
assign n2097____DOLLAR__5136 = oc8051_ROM_rdata_1[7:3] ;
assign n2098____DOLLAR__5142 =  { ( n2097____DOLLAR__5136 ) , ( 3'd0 ) }  ;
assign n2099____DOLLAR__5144 =  {3'd0 , n2097____DOLLAR__5136}  ;
assign n2100____DOLLAR__5146 =  ( n2099____DOLLAR__5144 ) + ( 8'd32 )  ;
assign n2101____DOLLAR__5147 =  ( n2096____DOLLAR__5134 ) ? ( n2098____DOLLAR__5142 ) : ( n2100____DOLLAR__5146 ) ;
assign n2102____DOLLAR__5150 =  ( n2101____DOLLAR__5147 ) == ( 8'd141 )  ;
assign n2103____DOLLAR__5155 = oc8051_ROM_rdata_1[7:7] ;
assign n2104____DOLLAR__5157 =  ( n2103____DOLLAR__5155 ) == ( 1'd1 )  ;
assign n2105____DOLLAR__5159 = oc8051_ROM_rdata_1[7:3] ;
assign n2106____DOLLAR__5165 =  { ( n2105____DOLLAR__5159 ) , ( 3'd0 ) }  ;
assign n2107____DOLLAR__5167 =  {3'd0 , n2105____DOLLAR__5159}  ;
assign n2108____DOLLAR__5169 =  ( n2107____DOLLAR__5167 ) + ( 8'd32 )  ;
assign n2109____DOLLAR__5170 =  ( n2104____DOLLAR__5157 ) ? ( n2106____DOLLAR__5165 ) : ( n2108____DOLLAR__5169 ) ;
assign n2110____DOLLAR__5173 =  ( n2109____DOLLAR__5170 ) == ( 8'd144 )  ;
assign n2111____DOLLAR__5178 = oc8051_ROM_rdata_1[7:7] ;
assign n2112____DOLLAR__5180 =  ( n2111____DOLLAR__5178 ) == ( 1'd1 )  ;
assign n2113____DOLLAR__5182 = oc8051_ROM_rdata_1[7:3] ;
assign n2114____DOLLAR__5188 =  { ( n2113____DOLLAR__5182 ) , ( 3'd0 ) }  ;
assign n2115____DOLLAR__5190 =  {3'd0 , n2113____DOLLAR__5182}  ;
assign n2116____DOLLAR__5192 =  ( n2115____DOLLAR__5190 ) + ( 8'd32 )  ;
assign n2117____DOLLAR__5193 =  ( n2112____DOLLAR__5180 ) ? ( n2114____DOLLAR__5188 ) : ( n2116____DOLLAR__5192 ) ;
assign n2118____DOLLAR__5196 =  ( n2117____DOLLAR__5193 ) == ( 8'd152 )  ;
assign n2119____DOLLAR__5201 = oc8051_ROM_rdata_1[7:7] ;
assign n2120____DOLLAR__5203 =  ( n2119____DOLLAR__5201 ) == ( 1'd1 )  ;
assign n2121____DOLLAR__5205 = oc8051_ROM_rdata_1[7:3] ;
assign n2122____DOLLAR__5211 =  { ( n2121____DOLLAR__5205 ) , ( 3'd0 ) }  ;
assign n2123____DOLLAR__5213 =  {3'd0 , n2121____DOLLAR__5205}  ;
assign n2124____DOLLAR__5215 =  ( n2123____DOLLAR__5213 ) + ( 8'd32 )  ;
assign n2125____DOLLAR__5216 =  ( n2120____DOLLAR__5203 ) ? ( n2122____DOLLAR__5211 ) : ( n2124____DOLLAR__5215 ) ;
assign n2126____DOLLAR__5219 =  ( n2125____DOLLAR__5216 ) == ( 8'd153 )  ;
assign n2127____DOLLAR__5224 = oc8051_ROM_rdata_1[7:7] ;
assign n2128____DOLLAR__5226 =  ( n2127____DOLLAR__5224 ) == ( 1'd1 )  ;
assign n2129____DOLLAR__5228 = oc8051_ROM_rdata_1[7:3] ;
assign n2130____DOLLAR__5234 =  { ( n2129____DOLLAR__5228 ) , ( 3'd0 ) }  ;
assign n2131____DOLLAR__5236 =  {3'd0 , n2129____DOLLAR__5228}  ;
assign n2132____DOLLAR__5238 =  ( n2131____DOLLAR__5236 ) + ( 8'd32 )  ;
assign n2133____DOLLAR__5239 =  ( n2128____DOLLAR__5226 ) ? ( n2130____DOLLAR__5234 ) : ( n2132____DOLLAR__5238 ) ;
assign n2134____DOLLAR__5242 =  ( n2133____DOLLAR__5239 ) == ( 8'd160 )  ;
assign n2135____DOLLAR__5247 = oc8051_ROM_rdata_1[7:7] ;
assign n2136____DOLLAR__5249 =  ( n2135____DOLLAR__5247 ) == ( 1'd1 )  ;
assign n2137____DOLLAR__5251 = oc8051_ROM_rdata_1[7:3] ;
assign n2138____DOLLAR__5257 =  { ( n2137____DOLLAR__5251 ) , ( 3'd0 ) }  ;
assign n2139____DOLLAR__5259 =  {3'd0 , n2137____DOLLAR__5251}  ;
assign n2140____DOLLAR__5261 =  ( n2139____DOLLAR__5259 ) + ( 8'd32 )  ;
assign n2141____DOLLAR__5262 =  ( n2136____DOLLAR__5249 ) ? ( n2138____DOLLAR__5257 ) : ( n2140____DOLLAR__5261 ) ;
assign n2142____DOLLAR__5265 =  ( n2141____DOLLAR__5262 ) == ( 8'd168 )  ;
assign n2143____DOLLAR__5270 = oc8051_ROM_rdata_1[7:7] ;
assign n2144____DOLLAR__5272 =  ( n2143____DOLLAR__5270 ) == ( 1'd1 )  ;
assign n2145____DOLLAR__5274 = oc8051_ROM_rdata_1[7:3] ;
assign n2146____DOLLAR__5280 =  { ( n2145____DOLLAR__5274 ) , ( 3'd0 ) }  ;
assign n2147____DOLLAR__5282 =  {3'd0 , n2145____DOLLAR__5274}  ;
assign n2148____DOLLAR__5284 =  ( n2147____DOLLAR__5282 ) + ( 8'd32 )  ;
assign n2149____DOLLAR__5285 =  ( n2144____DOLLAR__5272 ) ? ( n2146____DOLLAR__5280 ) : ( n2148____DOLLAR__5284 ) ;
assign n2150____DOLLAR__5288 =  ( n2149____DOLLAR__5285 ) == ( 8'd176 )  ;
assign n2151____DOLLAR__5293 = oc8051_ROM_rdata_1[7:7] ;
assign n2152____DOLLAR__5295 =  ( n2151____DOLLAR__5293 ) == ( 1'd1 )  ;
assign n2153____DOLLAR__5297 = oc8051_ROM_rdata_1[7:3] ;
assign n2154____DOLLAR__5303 =  { ( n2153____DOLLAR__5297 ) , ( 3'd0 ) }  ;
assign n2155____DOLLAR__5305 =  {3'd0 , n2153____DOLLAR__5297}  ;
assign n2156____DOLLAR__5307 =  ( n2155____DOLLAR__5305 ) + ( 8'd32 )  ;
assign n2157____DOLLAR__5308 =  ( n2152____DOLLAR__5295 ) ? ( n2154____DOLLAR__5303 ) : ( n2156____DOLLAR__5307 ) ;
assign n2158____DOLLAR__5311 =  ( n2157____DOLLAR__5308 ) == ( 8'd184 )  ;
assign n2159____DOLLAR__5316 = oc8051_ROM_rdata_1[7:7] ;
assign n2160____DOLLAR__5318 =  ( n2159____DOLLAR__5316 ) == ( 1'd1 )  ;
assign n2161____DOLLAR__5320 = oc8051_ROM_rdata_1[7:3] ;
assign n2162____DOLLAR__5326 =  { ( n2161____DOLLAR__5320 ) , ( 3'd0 ) }  ;
assign n2163____DOLLAR__5328 =  {3'd0 , n2161____DOLLAR__5320}  ;
assign n2164____DOLLAR__5330 =  ( n2163____DOLLAR__5328 ) + ( 8'd32 )  ;
assign n2165____DOLLAR__5331 =  ( n2160____DOLLAR__5318 ) ? ( n2162____DOLLAR__5326 ) : ( n2164____DOLLAR__5330 ) ;
assign n2166____DOLLAR__5334 =  ( n2165____DOLLAR__5331 ) == ( 8'd208 )  ;
assign n2167____DOLLAR__5339 = oc8051_ROM_rdata_1[7:7] ;
assign n2168____DOLLAR__5341 =  ( n2167____DOLLAR__5339 ) == ( 1'd1 )  ;
assign n2169____DOLLAR__5343 = oc8051_ROM_rdata_1[7:3] ;
assign n2170____DOLLAR__5349 =  { ( n2169____DOLLAR__5343 ) , ( 3'd0 ) }  ;
assign n2171____DOLLAR__5351 =  {3'd0 , n2169____DOLLAR__5343}  ;
assign n2172____DOLLAR__5353 =  ( n2171____DOLLAR__5351 ) + ( 8'd32 )  ;
assign n2173____DOLLAR__5354 =  ( n2168____DOLLAR__5341 ) ? ( n2170____DOLLAR__5349 ) : ( n2172____DOLLAR__5353 ) ;
assign n2174____DOLLAR__5357 =  ( n2173____DOLLAR__5354 ) == ( 8'd224 )  ;
assign n2175____DOLLAR__5362 = oc8051_ROM_rdata_1[7:7] ;
assign n2176____DOLLAR__5364 =  ( n2175____DOLLAR__5362 ) == ( 1'd1 )  ;
assign n2177____DOLLAR__5366 = oc8051_ROM_rdata_1[7:3] ;
assign n2178____DOLLAR__5372 =  { ( n2177____DOLLAR__5366 ) , ( 3'd0 ) }  ;
assign n2179____DOLLAR__5374 =  {3'd0 , n2177____DOLLAR__5366}  ;
assign n2180____DOLLAR__5376 =  ( n2179____DOLLAR__5374 ) + ( 8'd32 )  ;
assign n2181____DOLLAR__5377 =  ( n2176____DOLLAR__5364 ) ? ( n2178____DOLLAR__5372 ) : ( n2180____DOLLAR__5376 ) ;
assign n2182____DOLLAR__5380 =  ( n2181____DOLLAR__5377 ) == ( 8'd240 )  ;
assign n2183____DOLLAR__5384 =  ( n2182____DOLLAR__5380 ) ? ( B ) : ( 8'd0 ) ;
assign n2184____DOLLAR__5385 =  ( n2174____DOLLAR__5357 ) ? ( ACC ) : ( n2183____DOLLAR__5384 ) ;
assign n2185____DOLLAR__5386 =  ( n2166____DOLLAR__5334 ) ? ( PSW ) : ( n2184____DOLLAR__5385 ) ;
assign n2186____DOLLAR__5387 =  ( n2158____DOLLAR__5311 ) ? ( IP ) : ( n2185____DOLLAR__5386 ) ;
assign n2187____DOLLAR__5388 =  ( n2150____DOLLAR__5288 ) ? ( P3 ) : ( n2186____DOLLAR__5387 ) ;
assign n2188____DOLLAR__5389 =  ( n2142____DOLLAR__5265 ) ? ( IE ) : ( n2187____DOLLAR__5388 ) ;
assign n2189____DOLLAR__5390 =  ( n2134____DOLLAR__5242 ) ? ( P2 ) : ( n2188____DOLLAR__5389 ) ;
assign n2190____DOLLAR__5391 =  ( n2126____DOLLAR__5219 ) ? ( SBUF ) : ( n2189____DOLLAR__5390 ) ;
assign n2191____DOLLAR__5392 =  ( n2118____DOLLAR__5196 ) ? ( SCON ) : ( n2190____DOLLAR__5391 ) ;
assign n2192____DOLLAR__5393 =  ( n2110____DOLLAR__5173 ) ? ( P1 ) : ( n2191____DOLLAR__5392 ) ;
assign n2193____DOLLAR__5394 =  ( n2102____DOLLAR__5150 ) ? ( TH1 ) : ( n2192____DOLLAR__5393 ) ;
assign n2194____DOLLAR__5395 =  ( n2094____DOLLAR__5127 ) ? ( TL1 ) : ( n2193____DOLLAR__5394 ) ;
assign n2195____DOLLAR__5396 =  ( n2086____DOLLAR__5104 ) ? ( TH0 ) : ( n2194____DOLLAR__5395 ) ;
assign n2196____DOLLAR__5397 =  ( n2078____DOLLAR__5081 ) ? ( TL0 ) : ( n2195____DOLLAR__5396 ) ;
assign n2197____DOLLAR__5398 =  ( n2070____DOLLAR__5058 ) ? ( TMOD ) : ( n2196____DOLLAR__5397 ) ;
assign n2198____DOLLAR__5399 =  ( n2062____DOLLAR__5035 ) ? ( TCON ) : ( n2197____DOLLAR__5398 ) ;
assign n2199____DOLLAR__5400 =  ( n2054____DOLLAR__5012 ) ? ( PCON ) : ( n2198____DOLLAR__5399 ) ;
assign n2200____DOLLAR__5401 =  ( n2046____DOLLAR__4989 ) ? ( DPH ) : ( n2199____DOLLAR__5400 ) ;
assign n2201____DOLLAR__5402 =  ( n2038____DOLLAR__4966 ) ? ( DPL ) : ( n2200____DOLLAR__5401 ) ;
assign n2202____DOLLAR__5403 =  ( n2030____DOLLAR__4943 ) ? ( SP ) : ( n2201____DOLLAR__5402 ) ;
assign n2203____DOLLAR__5404 =  ( n2022____DOLLAR__4920 ) ? ( P0 ) : ( n2202____DOLLAR__5403 ) ;
assign n2204____DOLLAR__5405 =  ( n1973____DOLLAR__4868 ) ? ( n2014____DOLLAR__187168 ) : ( n2203____DOLLAR__5404 ) ;
assign n2205____DOLLAR__5406 =  ( n1964____DOLLAR__4844 ) & ( n2204____DOLLAR__5405 )  ;
assign n2206____DOLLAR__5407 = PSW[7:7] ;
assign n2207____DOLLAR__5409 =  {7'd0 , n2206____DOLLAR__5407}  ;
assign n2208____DOLLAR__5414 = oc8051_ROM_rdata_1[2:0] ;
assign n2209____DOLLAR__5416 =  {5'd0 , n2208____DOLLAR__5414}  ;
assign n2210____DOLLAR__5418 =  ( n2207____DOLLAR__5409 ) << ( n2209____DOLLAR__5416 )  ;
assign n2211____DOLLAR__5419 =  ( n2205____DOLLAR__5406 ) | ( n2210____DOLLAR__5418 )  ;
assign n2212____DOLLAR__5420 =  ( n1960____DOLLAR__4832 ) ? ( n2211____DOLLAR__5419 ) : ( SP ) ;
assign n2213____DOLLAR__5421 =  ( n1952____DOLLAR__4802 ) ? ( n2212____DOLLAR__5420 ) : ( SP ) ;
assign n2214____DOLLAR__5426 =  ( oc8051_ROM_rdata_0 ) == ( 8'd243 )  ;
assign n2215____DOLLAR__5430 =  ( oc8051_ROM_rdata_0 ) == ( 8'd227 )  ;
assign n2216____DOLLAR__5432 =  ( n2214____DOLLAR__5426 ) | ( n2215____DOLLAR__5430 )  ;
assign n2217____DOLLAR__5437 = PSW[4:3] ;
assign n2218____DOLLAR__5445 =  { ( n2217____DOLLAR__5437 ) , ( 3'd1 ) }  ;
assign n2219____DOLLAR__5451 =  { ( 3'd0 ) , ( n2218____DOLLAR__5445 ) }  ;
assign n2220____DOLLAR__192041 = n2219____DOLLAR__5451[3:0] ;
assign n2221____DOLLAR__192122 =  ( n2220____DOLLAR__192041 ) == ( 4'd15 )  ;
assign n2222____DOLLAR__192117 =  ( n2220____DOLLAR__192041 ) == ( 4'd14 )  ;
assign n2223____DOLLAR__192112 =  ( n2220____DOLLAR__192041 ) == ( 4'd13 )  ;
assign n2224____DOLLAR__192107 =  ( n2220____DOLLAR__192041 ) == ( 4'd12 )  ;
assign n2225____DOLLAR__192102 =  ( n2220____DOLLAR__192041 ) == ( 4'd11 )  ;
assign n2226____DOLLAR__192097 =  ( n2220____DOLLAR__192041 ) == ( 4'd10 )  ;
assign n2227____DOLLAR__192092 =  ( n2220____DOLLAR__192041 ) == ( 4'd9 )  ;
assign n2228____DOLLAR__192087 =  ( n2220____DOLLAR__192041 ) == ( 4'd8 )  ;
assign n2229____DOLLAR__192082 =  ( n2220____DOLLAR__192041 ) == ( 4'd7 )  ;
assign n2230____DOLLAR__192077 =  ( n2220____DOLLAR__192041 ) == ( 4'd6 )  ;
assign n2231____DOLLAR__192072 =  ( n2220____DOLLAR__192041 ) == ( 4'd5 )  ;
assign n2232____DOLLAR__192067 =  ( n2220____DOLLAR__192041 ) == ( 4'd4 )  ;
assign n2233____DOLLAR__192062 =  ( n2220____DOLLAR__192041 ) == ( 4'd3 )  ;
assign n2234____DOLLAR__192057 =  ( n2220____DOLLAR__192041 ) == ( 4'd2 )  ;
assign n2235____DOLLAR__192052 =  ( n2220____DOLLAR__192041 ) == ( 4'd1 )  ;
assign n2236____DOLLAR__192047 =  ( n2220____DOLLAR__192041 ) == ( 4'd0 )  ;
assign n2237____DOLLAR__192049 =  ( n2236____DOLLAR__192047 ) ? ( oc8051_IRAM_data_0 ) : ( 8'd0 ) ;
assign n2238____DOLLAR__192054 =  ( n2235____DOLLAR__192052 ) ? ( oc8051_IRAM_data_1 ) : ( n2237____DOLLAR__192049 ) ;
assign n2239____DOLLAR__192059 =  ( n2234____DOLLAR__192057 ) ? ( oc8051_IRAM_data_2 ) : ( n2238____DOLLAR__192054 ) ;
assign n2240____DOLLAR__192064 =  ( n2233____DOLLAR__192062 ) ? ( oc8051_IRAM_data_3 ) : ( n2239____DOLLAR__192059 ) ;
assign n2241____DOLLAR__192069 =  ( n2232____DOLLAR__192067 ) ? ( oc8051_IRAM_data_4 ) : ( n2240____DOLLAR__192064 ) ;
assign n2242____DOLLAR__192074 =  ( n2231____DOLLAR__192072 ) ? ( oc8051_IRAM_data_5 ) : ( n2241____DOLLAR__192069 ) ;
assign n2243____DOLLAR__192079 =  ( n2230____DOLLAR__192077 ) ? ( oc8051_IRAM_data_6 ) : ( n2242____DOLLAR__192074 ) ;
assign n2244____DOLLAR__192084 =  ( n2229____DOLLAR__192082 ) ? ( oc8051_IRAM_data_7 ) : ( n2243____DOLLAR__192079 ) ;
assign n2245____DOLLAR__192089 =  ( n2228____DOLLAR__192087 ) ? ( oc8051_IRAM_data_8 ) : ( n2244____DOLLAR__192084 ) ;
assign n2246____DOLLAR__192094 =  ( n2227____DOLLAR__192092 ) ? ( oc8051_IRAM_data_9 ) : ( n2245____DOLLAR__192089 ) ;
assign n2247____DOLLAR__192099 =  ( n2226____DOLLAR__192097 ) ? ( oc8051_IRAM_data_10 ) : ( n2246____DOLLAR__192094 ) ;
assign n2248____DOLLAR__192104 =  ( n2225____DOLLAR__192102 ) ? ( oc8051_IRAM_data_11 ) : ( n2247____DOLLAR__192099 ) ;
assign n2249____DOLLAR__192109 =  ( n2224____DOLLAR__192107 ) ? ( oc8051_IRAM_data_12 ) : ( n2248____DOLLAR__192104 ) ;
assign n2250____DOLLAR__192114 =  ( n2223____DOLLAR__192112 ) ? ( oc8051_IRAM_data_13 ) : ( n2249____DOLLAR__192109 ) ;
assign n2251____DOLLAR__192119 =  ( n2222____DOLLAR__192117 ) ? ( oc8051_IRAM_data_14 ) : ( n2250____DOLLAR__192114 ) ;
assign n2252____DOLLAR__192124 =  ( n2221____DOLLAR__192122 ) ? ( oc8051_IRAM_data_15 ) : ( n2251____DOLLAR__192119 ) ;
assign n2253____DOLLAR__5459 =  { ( 8'd0 ) , ( n2252____DOLLAR__192124 ) }  ;
assign n2254____DOLLAR__5465 =  ( oc8051_ROM_rdata_0 ) == ( 8'd242 )  ;
assign n2255____DOLLAR__5469 =  ( oc8051_ROM_rdata_0 ) == ( 8'd226 )  ;
assign n2256____DOLLAR__5471 =  ( n2254____DOLLAR__5465 ) | ( n2255____DOLLAR__5469 )  ;
assign n2257____DOLLAR__5476 = PSW[4:3] ;
assign n2258____DOLLAR__5484 =  { ( n2257____DOLLAR__5476 ) , ( 3'd0 ) }  ;
assign n2259____DOLLAR__5490 =  { ( 3'd0 ) , ( n2258____DOLLAR__5484 ) }  ;
assign n2260____DOLLAR__192149 = n2259____DOLLAR__5490[3:0] ;
assign n2261____DOLLAR__192230 =  ( n2260____DOLLAR__192149 ) == ( 4'd15 )  ;
assign n2262____DOLLAR__192225 =  ( n2260____DOLLAR__192149 ) == ( 4'd14 )  ;
assign n2263____DOLLAR__192220 =  ( n2260____DOLLAR__192149 ) == ( 4'd13 )  ;
assign n2264____DOLLAR__192215 =  ( n2260____DOLLAR__192149 ) == ( 4'd12 )  ;
assign n2265____DOLLAR__192210 =  ( n2260____DOLLAR__192149 ) == ( 4'd11 )  ;
assign n2266____DOLLAR__192205 =  ( n2260____DOLLAR__192149 ) == ( 4'd10 )  ;
assign n2267____DOLLAR__192200 =  ( n2260____DOLLAR__192149 ) == ( 4'd9 )  ;
assign n2268____DOLLAR__192195 =  ( n2260____DOLLAR__192149 ) == ( 4'd8 )  ;
assign n2269____DOLLAR__192190 =  ( n2260____DOLLAR__192149 ) == ( 4'd7 )  ;
assign n2270____DOLLAR__192185 =  ( n2260____DOLLAR__192149 ) == ( 4'd6 )  ;
assign n2271____DOLLAR__192180 =  ( n2260____DOLLAR__192149 ) == ( 4'd5 )  ;
assign n2272____DOLLAR__192175 =  ( n2260____DOLLAR__192149 ) == ( 4'd4 )  ;
assign n2273____DOLLAR__192170 =  ( n2260____DOLLAR__192149 ) == ( 4'd3 )  ;
assign n2274____DOLLAR__192165 =  ( n2260____DOLLAR__192149 ) == ( 4'd2 )  ;
assign n2275____DOLLAR__192160 =  ( n2260____DOLLAR__192149 ) == ( 4'd1 )  ;
assign n2276____DOLLAR__192155 =  ( n2260____DOLLAR__192149 ) == ( 4'd0 )  ;
assign n2277____DOLLAR__192157 =  ( n2276____DOLLAR__192155 ) ? ( oc8051_IRAM_data_0 ) : ( 8'd0 ) ;
assign n2278____DOLLAR__192162 =  ( n2275____DOLLAR__192160 ) ? ( oc8051_IRAM_data_1 ) : ( n2277____DOLLAR__192157 ) ;
assign n2279____DOLLAR__192167 =  ( n2274____DOLLAR__192165 ) ? ( oc8051_IRAM_data_2 ) : ( n2278____DOLLAR__192162 ) ;
assign n2280____DOLLAR__192172 =  ( n2273____DOLLAR__192170 ) ? ( oc8051_IRAM_data_3 ) : ( n2279____DOLLAR__192167 ) ;
assign n2281____DOLLAR__192177 =  ( n2272____DOLLAR__192175 ) ? ( oc8051_IRAM_data_4 ) : ( n2280____DOLLAR__192172 ) ;
assign n2282____DOLLAR__192182 =  ( n2271____DOLLAR__192180 ) ? ( oc8051_IRAM_data_5 ) : ( n2281____DOLLAR__192177 ) ;
assign n2283____DOLLAR__192187 =  ( n2270____DOLLAR__192185 ) ? ( oc8051_IRAM_data_6 ) : ( n2282____DOLLAR__192182 ) ;
assign n2284____DOLLAR__192192 =  ( n2269____DOLLAR__192190 ) ? ( oc8051_IRAM_data_7 ) : ( n2283____DOLLAR__192187 ) ;
assign n2285____DOLLAR__192197 =  ( n2268____DOLLAR__192195 ) ? ( oc8051_IRAM_data_8 ) : ( n2284____DOLLAR__192192 ) ;
assign n2286____DOLLAR__192202 =  ( n2267____DOLLAR__192200 ) ? ( oc8051_IRAM_data_9 ) : ( n2285____DOLLAR__192197 ) ;
assign n2287____DOLLAR__192207 =  ( n2266____DOLLAR__192205 ) ? ( oc8051_IRAM_data_10 ) : ( n2286____DOLLAR__192202 ) ;
assign n2288____DOLLAR__192212 =  ( n2265____DOLLAR__192210 ) ? ( oc8051_IRAM_data_11 ) : ( n2287____DOLLAR__192207 ) ;
assign n2289____DOLLAR__192217 =  ( n2264____DOLLAR__192215 ) ? ( oc8051_IRAM_data_12 ) : ( n2288____DOLLAR__192212 ) ;
assign n2290____DOLLAR__192222 =  ( n2263____DOLLAR__192220 ) ? ( oc8051_IRAM_data_13 ) : ( n2289____DOLLAR__192217 ) ;
assign n2291____DOLLAR__192227 =  ( n2262____DOLLAR__192225 ) ? ( oc8051_IRAM_data_14 ) : ( n2290____DOLLAR__192222 ) ;
assign n2292____DOLLAR__192232 =  ( n2261____DOLLAR__192230 ) ? ( oc8051_IRAM_data_15 ) : ( n2291____DOLLAR__192227 ) ;
assign n2293____DOLLAR__5498 =  { ( 8'd0 ) , ( n2292____DOLLAR__192232 ) }  ;
assign n2294____DOLLAR__5504 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign n2295____DOLLAR__5508 =  ( oc8051_ROM_rdata_0 ) == ( 8'd224 )  ;
assign n2296____DOLLAR__5510 =  ( n2294____DOLLAR__5504 ) | ( n2295____DOLLAR__5508 )  ;
assign n2297____DOLLAR__5515 =  { ( DPH ) , ( DPL ) }  ;
assign n2298____DOLLAR__5521 =  ( oc8051_ROM_rdata_0 ) == ( 8'd255 )  ;
assign n2299____DOLLAR__5525 =  ( oc8051_ROM_rdata_0 ) == ( 8'd254 )  ;
assign n2300____DOLLAR__5529 =  ( oc8051_ROM_rdata_0 ) == ( 8'd253 )  ;
assign n2301____DOLLAR__5533 =  ( oc8051_ROM_rdata_0 ) == ( 8'd252 )  ;
assign n2302____DOLLAR__5537 =  ( oc8051_ROM_rdata_0 ) == ( 8'd251 )  ;
assign n2303____DOLLAR__5541 =  ( oc8051_ROM_rdata_0 ) == ( 8'd250 )  ;
assign n2304____DOLLAR__5545 =  ( oc8051_ROM_rdata_0 ) == ( 8'd249 )  ;
assign n2305____DOLLAR__5549 =  ( oc8051_ROM_rdata_0 ) == ( 8'd248 )  ;
assign n2306____DOLLAR__5553 =  ( oc8051_ROM_rdata_0 ) == ( 8'd247 )  ;
assign n2307____DOLLAR__5557 =  ( oc8051_ROM_rdata_0 ) == ( 8'd246 )  ;
assign n2308____DOLLAR__5561 =  ( oc8051_ROM_rdata_0 ) == ( 8'd245 )  ;
assign n2309____DOLLAR__5565 =  ( oc8051_ROM_rdata_0 ) == ( 8'd244 )  ;
assign n2310____DOLLAR__5569 =  ( oc8051_ROM_rdata_0 ) == ( 8'd241 )  ;
assign n2311____DOLLAR__5573 =  ( oc8051_ROM_rdata_0 ) == ( 8'd239 )  ;
assign n2312____DOLLAR__5577 =  ( oc8051_ROM_rdata_0 ) == ( 8'd238 )  ;
assign n2313____DOLLAR__5581 =  ( oc8051_ROM_rdata_0 ) == ( 8'd237 )  ;
assign n2314____DOLLAR__5585 =  ( oc8051_ROM_rdata_0 ) == ( 8'd236 )  ;
assign n2315____DOLLAR__5589 =  ( oc8051_ROM_rdata_0 ) == ( 8'd235 )  ;
assign n2316____DOLLAR__5593 =  ( oc8051_ROM_rdata_0 ) == ( 8'd234 )  ;
assign n2317____DOLLAR__5597 =  ( oc8051_ROM_rdata_0 ) == ( 8'd233 )  ;
assign n2318____DOLLAR__5601 =  ( oc8051_ROM_rdata_0 ) == ( 8'd232 )  ;
assign n2319____DOLLAR__5605 =  ( oc8051_ROM_rdata_0 ) == ( 8'd231 )  ;
assign n2320____DOLLAR__5609 =  ( oc8051_ROM_rdata_0 ) == ( 8'd230 )  ;
assign n2321____DOLLAR__5613 =  ( oc8051_ROM_rdata_0 ) == ( 8'd229 )  ;
assign n2322____DOLLAR__5617 =  ( oc8051_ROM_rdata_0 ) == ( 8'd228 )  ;
assign n2323____DOLLAR__5621 =  ( oc8051_ROM_rdata_0 ) == ( 8'd225 )  ;
assign n2324____DOLLAR__5625 =  ( oc8051_ROM_rdata_0 ) == ( 8'd223 )  ;
assign n2325____DOLLAR__5629 =  ( oc8051_ROM_rdata_0 ) == ( 8'd222 )  ;
assign n2326____DOLLAR__5633 =  ( oc8051_ROM_rdata_0 ) == ( 8'd221 )  ;
assign n2327____DOLLAR__5637 =  ( oc8051_ROM_rdata_0 ) == ( 8'd220 )  ;
assign n2328____DOLLAR__5641 =  ( oc8051_ROM_rdata_0 ) == ( 8'd219 )  ;
assign n2329____DOLLAR__5645 =  ( oc8051_ROM_rdata_0 ) == ( 8'd218 )  ;
assign n2330____DOLLAR__5649 =  ( oc8051_ROM_rdata_0 ) == ( 8'd217 )  ;
assign n2331____DOLLAR__5653 =  ( oc8051_ROM_rdata_0 ) == ( 8'd216 )  ;
assign n2332____DOLLAR__5657 =  ( oc8051_ROM_rdata_0 ) == ( 8'd215 )  ;
assign n2333____DOLLAR__5661 =  ( oc8051_ROM_rdata_0 ) == ( 8'd214 )  ;
assign n2334____DOLLAR__5665 =  ( oc8051_ROM_rdata_0 ) == ( 8'd213 )  ;
assign n2335____DOLLAR__5669 =  ( oc8051_ROM_rdata_0 ) == ( 8'd212 )  ;
assign n2336____DOLLAR__5673 =  ( oc8051_ROM_rdata_0 ) == ( 8'd211 )  ;
assign n2337____DOLLAR__5677 =  ( oc8051_ROM_rdata_0 ) == ( 8'd210 )  ;
assign n2338____DOLLAR__5681 =  ( oc8051_ROM_rdata_0 ) == ( 8'd209 )  ;
assign n2339____DOLLAR__5685 =  ( oc8051_ROM_rdata_0 ) == ( 8'd208 )  ;
assign n2340____DOLLAR__5689 =  ( oc8051_ROM_rdata_0 ) == ( 8'd207 )  ;
assign n2341____DOLLAR__5693 =  ( oc8051_ROM_rdata_0 ) == ( 8'd206 )  ;
assign n2342____DOLLAR__5697 =  ( oc8051_ROM_rdata_0 ) == ( 8'd205 )  ;
assign n2343____DOLLAR__5701 =  ( oc8051_ROM_rdata_0 ) == ( 8'd204 )  ;
assign n2344____DOLLAR__5705 =  ( oc8051_ROM_rdata_0 ) == ( 8'd203 )  ;
assign n2345____DOLLAR__5709 =  ( oc8051_ROM_rdata_0 ) == ( 8'd202 )  ;
assign n2346____DOLLAR__5713 =  ( oc8051_ROM_rdata_0 ) == ( 8'd201 )  ;
assign n2347____DOLLAR__5717 =  ( oc8051_ROM_rdata_0 ) == ( 8'd200 )  ;
assign n2348____DOLLAR__5721 =  ( oc8051_ROM_rdata_0 ) == ( 8'd199 )  ;
assign n2349____DOLLAR__5725 =  ( oc8051_ROM_rdata_0 ) == ( 8'd198 )  ;
assign n2350____DOLLAR__5729 =  ( oc8051_ROM_rdata_0 ) == ( 8'd197 )  ;
assign n2351____DOLLAR__5733 =  ( oc8051_ROM_rdata_0 ) == ( 8'd196 )  ;
assign n2352____DOLLAR__5737 =  ( oc8051_ROM_rdata_0 ) == ( 8'd195 )  ;
assign n2353____DOLLAR__5741 =  ( oc8051_ROM_rdata_0 ) == ( 8'd194 )  ;
assign n2354____DOLLAR__5745 =  ( oc8051_ROM_rdata_0 ) == ( 8'd193 )  ;
assign n2355____DOLLAR__5749 =  ( oc8051_ROM_rdata_0 ) == ( 8'd192 )  ;
assign n2356____DOLLAR__5753 =  ( oc8051_ROM_rdata_0 ) == ( 8'd191 )  ;
assign n2357____DOLLAR__5757 =  ( oc8051_ROM_rdata_0 ) == ( 8'd190 )  ;
assign n2358____DOLLAR__5761 =  ( oc8051_ROM_rdata_0 ) == ( 8'd189 )  ;
assign n2359____DOLLAR__5765 =  ( oc8051_ROM_rdata_0 ) == ( 8'd188 )  ;
assign n2360____DOLLAR__5769 =  ( oc8051_ROM_rdata_0 ) == ( 8'd187 )  ;
assign n2361____DOLLAR__5773 =  ( oc8051_ROM_rdata_0 ) == ( 8'd186 )  ;
assign n2362____DOLLAR__5777 =  ( oc8051_ROM_rdata_0 ) == ( 8'd185 )  ;
assign n2363____DOLLAR__5781 =  ( oc8051_ROM_rdata_0 ) == ( 8'd184 )  ;
assign n2364____DOLLAR__5785 =  ( oc8051_ROM_rdata_0 ) == ( 8'd183 )  ;
assign n2365____DOLLAR__5789 =  ( oc8051_ROM_rdata_0 ) == ( 8'd182 )  ;
assign n2366____DOLLAR__5793 =  ( oc8051_ROM_rdata_0 ) == ( 8'd181 )  ;
assign n2367____DOLLAR__5797 =  ( oc8051_ROM_rdata_0 ) == ( 8'd180 )  ;
assign n2368____DOLLAR__5801 =  ( oc8051_ROM_rdata_0 ) == ( 8'd179 )  ;
assign n2369____DOLLAR__5805 =  ( oc8051_ROM_rdata_0 ) == ( 8'd178 )  ;
assign n2370____DOLLAR__5809 =  ( oc8051_ROM_rdata_0 ) == ( 8'd177 )  ;
assign n2371____DOLLAR__5813 =  ( oc8051_ROM_rdata_0 ) == ( 8'd176 )  ;
assign n2372____DOLLAR__5817 =  ( oc8051_ROM_rdata_0 ) == ( 8'd175 )  ;
assign n2373____DOLLAR__5821 =  ( oc8051_ROM_rdata_0 ) == ( 8'd174 )  ;
assign n2374____DOLLAR__5825 =  ( oc8051_ROM_rdata_0 ) == ( 8'd173 )  ;
assign n2375____DOLLAR__5829 =  ( oc8051_ROM_rdata_0 ) == ( 8'd172 )  ;
assign n2376____DOLLAR__5833 =  ( oc8051_ROM_rdata_0 ) == ( 8'd171 )  ;
assign n2377____DOLLAR__5837 =  ( oc8051_ROM_rdata_0 ) == ( 8'd170 )  ;
assign n2378____DOLLAR__5841 =  ( oc8051_ROM_rdata_0 ) == ( 8'd169 )  ;
assign n2379____DOLLAR__5845 =  ( oc8051_ROM_rdata_0 ) == ( 8'd168 )  ;
assign n2380____DOLLAR__5849 =  ( oc8051_ROM_rdata_0 ) == ( 8'd167 )  ;
assign n2381____DOLLAR__5853 =  ( oc8051_ROM_rdata_0 ) == ( 8'd166 )  ;
assign n2382____DOLLAR__5857 =  ( oc8051_ROM_rdata_0 ) == ( 8'd165 )  ;
assign n2383____DOLLAR__5861 =  ( oc8051_ROM_rdata_0 ) == ( 8'd164 )  ;
assign n2384____DOLLAR__5865 =  ( oc8051_ROM_rdata_0 ) == ( 8'd163 )  ;
assign n2385____DOLLAR__5869 =  ( oc8051_ROM_rdata_0 ) == ( 8'd162 )  ;
assign n2386____DOLLAR__5873 =  ( oc8051_ROM_rdata_0 ) == ( 8'd161 )  ;
assign n2387____DOLLAR__5877 =  ( oc8051_ROM_rdata_0 ) == ( 8'd160 )  ;
assign n2388____DOLLAR__5881 =  ( oc8051_ROM_rdata_0 ) == ( 8'd159 )  ;
assign n2389____DOLLAR__5885 =  ( oc8051_ROM_rdata_0 ) == ( 8'd158 )  ;
assign n2390____DOLLAR__5889 =  ( oc8051_ROM_rdata_0 ) == ( 8'd157 )  ;
assign n2391____DOLLAR__5893 =  ( oc8051_ROM_rdata_0 ) == ( 8'd156 )  ;
assign n2392____DOLLAR__5897 =  ( oc8051_ROM_rdata_0 ) == ( 8'd155 )  ;
assign n2393____DOLLAR__5901 =  ( oc8051_ROM_rdata_0 ) == ( 8'd154 )  ;
assign n2394____DOLLAR__5905 =  ( oc8051_ROM_rdata_0 ) == ( 8'd153 )  ;
assign n2395____DOLLAR__5909 =  ( oc8051_ROM_rdata_0 ) == ( 8'd152 )  ;
assign n2396____DOLLAR__5913 =  ( oc8051_ROM_rdata_0 ) == ( 8'd151 )  ;
assign n2397____DOLLAR__5917 =  ( oc8051_ROM_rdata_0 ) == ( 8'd150 )  ;
assign n2398____DOLLAR__5921 =  ( oc8051_ROM_rdata_0 ) == ( 8'd149 )  ;
assign n2399____DOLLAR__5925 =  ( oc8051_ROM_rdata_0 ) == ( 8'd148 )  ;
assign n2400____DOLLAR__5929 =  ( oc8051_ROM_rdata_0 ) == ( 8'd147 )  ;
assign n2401____DOLLAR__5933 =  ( oc8051_ROM_rdata_0 ) == ( 8'd146 )  ;
assign n2402____DOLLAR__5937 =  ( oc8051_ROM_rdata_0 ) == ( 8'd145 )  ;
assign n2403____DOLLAR__5941 =  ( oc8051_ROM_rdata_0 ) == ( 8'd144 )  ;
assign n2404____DOLLAR__5945 =  ( oc8051_ROM_rdata_0 ) == ( 8'd143 )  ;
assign n2405____DOLLAR__5949 =  ( oc8051_ROM_rdata_0 ) == ( 8'd142 )  ;
assign n2406____DOLLAR__5953 =  ( oc8051_ROM_rdata_0 ) == ( 8'd141 )  ;
assign n2407____DOLLAR__5957 =  ( oc8051_ROM_rdata_0 ) == ( 8'd140 )  ;
assign n2408____DOLLAR__5961 =  ( oc8051_ROM_rdata_0 ) == ( 8'd139 )  ;
assign n2409____DOLLAR__5965 =  ( oc8051_ROM_rdata_0 ) == ( 8'd138 )  ;
assign n2410____DOLLAR__5969 =  ( oc8051_ROM_rdata_0 ) == ( 8'd137 )  ;
assign n2411____DOLLAR__5973 =  ( oc8051_ROM_rdata_0 ) == ( 8'd136 )  ;
assign n2412____DOLLAR__5977 =  ( oc8051_ROM_rdata_0 ) == ( 8'd135 )  ;
assign n2413____DOLLAR__5981 =  ( oc8051_ROM_rdata_0 ) == ( 8'd134 )  ;
assign n2414____DOLLAR__5985 =  ( oc8051_ROM_rdata_0 ) == ( 8'd133 )  ;
assign n2415____DOLLAR__5989 =  ( oc8051_ROM_rdata_0 ) == ( 8'd132 )  ;
assign n2416____DOLLAR__5993 =  ( oc8051_ROM_rdata_0 ) == ( 8'd131 )  ;
assign n2417____DOLLAR__5997 =  ( oc8051_ROM_rdata_0 ) == ( 8'd130 )  ;
assign n2418____DOLLAR__6001 =  ( oc8051_ROM_rdata_0 ) == ( 8'd129 )  ;
assign n2419____DOLLAR__6005 =  ( oc8051_ROM_rdata_0 ) == ( 8'd128 )  ;
assign n2420____DOLLAR__6009 =  ( oc8051_ROM_rdata_0 ) == ( 8'd127 )  ;
assign n2421____DOLLAR__6013 =  ( oc8051_ROM_rdata_0 ) == ( 8'd126 )  ;
assign n2422____DOLLAR__6017 =  ( oc8051_ROM_rdata_0 ) == ( 8'd125 )  ;
assign n2423____DOLLAR__6021 =  ( oc8051_ROM_rdata_0 ) == ( 8'd124 )  ;
assign n2424____DOLLAR__6025 =  ( oc8051_ROM_rdata_0 ) == ( 8'd123 )  ;
assign n2425____DOLLAR__6029 =  ( oc8051_ROM_rdata_0 ) == ( 8'd122 )  ;
assign n2426____DOLLAR__6033 =  ( oc8051_ROM_rdata_0 ) == ( 8'd121 )  ;
assign n2427____DOLLAR__6037 =  ( oc8051_ROM_rdata_0 ) == ( 8'd120 )  ;
assign n2428____DOLLAR__6041 =  ( oc8051_ROM_rdata_0 ) == ( 8'd119 )  ;
assign n2429____DOLLAR__6045 =  ( oc8051_ROM_rdata_0 ) == ( 8'd118 )  ;
assign n2430____DOLLAR__6049 =  ( oc8051_ROM_rdata_0 ) == ( 8'd117 )  ;
assign n2431____DOLLAR__6053 =  ( oc8051_ROM_rdata_0 ) == ( 8'd116 )  ;
assign n2432____DOLLAR__6057 =  ( oc8051_ROM_rdata_0 ) == ( 8'd115 )  ;
assign n2433____DOLLAR__6061 =  ( oc8051_ROM_rdata_0 ) == ( 8'd114 )  ;
assign n2434____DOLLAR__6065 =  ( oc8051_ROM_rdata_0 ) == ( 8'd113 )  ;
assign n2435____DOLLAR__6069 =  ( oc8051_ROM_rdata_0 ) == ( 8'd112 )  ;
assign n2436____DOLLAR__6073 =  ( oc8051_ROM_rdata_0 ) == ( 8'd111 )  ;
assign n2437____DOLLAR__6077 =  ( oc8051_ROM_rdata_0 ) == ( 8'd110 )  ;
assign n2438____DOLLAR__6081 =  ( oc8051_ROM_rdata_0 ) == ( 8'd109 )  ;
assign n2439____DOLLAR__6085 =  ( oc8051_ROM_rdata_0 ) == ( 8'd108 )  ;
assign n2440____DOLLAR__6089 =  ( oc8051_ROM_rdata_0 ) == ( 8'd107 )  ;
assign n2441____DOLLAR__6093 =  ( oc8051_ROM_rdata_0 ) == ( 8'd106 )  ;
assign n2442____DOLLAR__6097 =  ( oc8051_ROM_rdata_0 ) == ( 8'd105 )  ;
assign n2443____DOLLAR__6101 =  ( oc8051_ROM_rdata_0 ) == ( 8'd104 )  ;
assign n2444____DOLLAR__6105 =  ( oc8051_ROM_rdata_0 ) == ( 8'd103 )  ;
assign n2445____DOLLAR__6109 =  ( oc8051_ROM_rdata_0 ) == ( 8'd102 )  ;
assign n2446____DOLLAR__6113 =  ( oc8051_ROM_rdata_0 ) == ( 8'd101 )  ;
assign n2447____DOLLAR__6117 =  ( oc8051_ROM_rdata_0 ) == ( 8'd100 )  ;
assign n2448____DOLLAR__6121 =  ( oc8051_ROM_rdata_0 ) == ( 8'd99 )  ;
assign n2449____DOLLAR__6125 =  ( oc8051_ROM_rdata_0 ) == ( 8'd98 )  ;
assign n2450____DOLLAR__6129 =  ( oc8051_ROM_rdata_0 ) == ( 8'd97 )  ;
assign n2451____DOLLAR__6133 =  ( oc8051_ROM_rdata_0 ) == ( 8'd96 )  ;
assign n2452____DOLLAR__6137 =  ( oc8051_ROM_rdata_0 ) == ( 8'd95 )  ;
assign n2453____DOLLAR__6141 =  ( oc8051_ROM_rdata_0 ) == ( 8'd94 )  ;
assign n2454____DOLLAR__6145 =  ( oc8051_ROM_rdata_0 ) == ( 8'd93 )  ;
assign n2455____DOLLAR__6149 =  ( oc8051_ROM_rdata_0 ) == ( 8'd92 )  ;
assign n2456____DOLLAR__6153 =  ( oc8051_ROM_rdata_0 ) == ( 8'd91 )  ;
assign n2457____DOLLAR__6157 =  ( oc8051_ROM_rdata_0 ) == ( 8'd90 )  ;
assign n2458____DOLLAR__6161 =  ( oc8051_ROM_rdata_0 ) == ( 8'd89 )  ;
assign n2459____DOLLAR__6165 =  ( oc8051_ROM_rdata_0 ) == ( 8'd88 )  ;
assign n2460____DOLLAR__6169 =  ( oc8051_ROM_rdata_0 ) == ( 8'd87 )  ;
assign n2461____DOLLAR__6173 =  ( oc8051_ROM_rdata_0 ) == ( 8'd86 )  ;
assign n2462____DOLLAR__6177 =  ( oc8051_ROM_rdata_0 ) == ( 8'd85 )  ;
assign n2463____DOLLAR__6181 =  ( oc8051_ROM_rdata_0 ) == ( 8'd84 )  ;
assign n2464____DOLLAR__6185 =  ( oc8051_ROM_rdata_0 ) == ( 8'd83 )  ;
assign n2465____DOLLAR__6189 =  ( oc8051_ROM_rdata_0 ) == ( 8'd82 )  ;
assign n2466____DOLLAR__6193 =  ( oc8051_ROM_rdata_0 ) == ( 8'd81 )  ;
assign n2467____DOLLAR__6197 =  ( oc8051_ROM_rdata_0 ) == ( 8'd80 )  ;
assign n2468____DOLLAR__6201 =  ( oc8051_ROM_rdata_0 ) == ( 8'd79 )  ;
assign n2469____DOLLAR__6205 =  ( oc8051_ROM_rdata_0 ) == ( 8'd78 )  ;
assign n2470____DOLLAR__6209 =  ( oc8051_ROM_rdata_0 ) == ( 8'd77 )  ;
assign n2471____DOLLAR__6213 =  ( oc8051_ROM_rdata_0 ) == ( 8'd76 )  ;
assign n2472____DOLLAR__6217 =  ( oc8051_ROM_rdata_0 ) == ( 8'd75 )  ;
assign n2473____DOLLAR__6221 =  ( oc8051_ROM_rdata_0 ) == ( 8'd74 )  ;
assign n2474____DOLLAR__6225 =  ( oc8051_ROM_rdata_0 ) == ( 8'd73 )  ;
assign n2475____DOLLAR__6229 =  ( oc8051_ROM_rdata_0 ) == ( 8'd72 )  ;
assign n2476____DOLLAR__6233 =  ( oc8051_ROM_rdata_0 ) == ( 8'd71 )  ;
assign n2477____DOLLAR__6237 =  ( oc8051_ROM_rdata_0 ) == ( 8'd70 )  ;
assign n2478____DOLLAR__6241 =  ( oc8051_ROM_rdata_0 ) == ( 8'd69 )  ;
assign n2479____DOLLAR__6245 =  ( oc8051_ROM_rdata_0 ) == ( 8'd68 )  ;
assign n2480____DOLLAR__6249 =  ( oc8051_ROM_rdata_0 ) == ( 8'd67 )  ;
assign n2481____DOLLAR__6253 =  ( oc8051_ROM_rdata_0 ) == ( 8'd66 )  ;
assign n2482____DOLLAR__6257 =  ( oc8051_ROM_rdata_0 ) == ( 8'd65 )  ;
assign n2483____DOLLAR__6261 =  ( oc8051_ROM_rdata_0 ) == ( 8'd64 )  ;
assign n2484____DOLLAR__6265 =  ( oc8051_ROM_rdata_0 ) == ( 8'd63 )  ;
assign n2485____DOLLAR__6269 =  ( oc8051_ROM_rdata_0 ) == ( 8'd62 )  ;
assign n2486____DOLLAR__6273 =  ( oc8051_ROM_rdata_0 ) == ( 8'd61 )  ;
assign n2487____DOLLAR__6277 =  ( oc8051_ROM_rdata_0 ) == ( 8'd60 )  ;
assign n2488____DOLLAR__6281 =  ( oc8051_ROM_rdata_0 ) == ( 8'd59 )  ;
assign n2489____DOLLAR__6285 =  ( oc8051_ROM_rdata_0 ) == ( 8'd58 )  ;
assign n2490____DOLLAR__6289 =  ( oc8051_ROM_rdata_0 ) == ( 8'd57 )  ;
assign n2491____DOLLAR__6293 =  ( oc8051_ROM_rdata_0 ) == ( 8'd56 )  ;
assign n2492____DOLLAR__6297 =  ( oc8051_ROM_rdata_0 ) == ( 8'd55 )  ;
assign n2493____DOLLAR__6301 =  ( oc8051_ROM_rdata_0 ) == ( 8'd54 )  ;
assign n2494____DOLLAR__6305 =  ( oc8051_ROM_rdata_0 ) == ( 8'd53 )  ;
assign n2495____DOLLAR__6309 =  ( oc8051_ROM_rdata_0 ) == ( 8'd52 )  ;
assign n2496____DOLLAR__6313 =  ( oc8051_ROM_rdata_0 ) == ( 8'd51 )  ;
assign n2497____DOLLAR__6317 =  ( oc8051_ROM_rdata_0 ) == ( 8'd50 )  ;
assign n2498____DOLLAR__6321 =  ( oc8051_ROM_rdata_0 ) == ( 8'd49 )  ;
assign n2499____DOLLAR__6325 =  ( oc8051_ROM_rdata_0 ) == ( 8'd48 )  ;
assign n2500____DOLLAR__6329 =  ( oc8051_ROM_rdata_0 ) == ( 8'd47 )  ;
assign n2501____DOLLAR__6333 =  ( oc8051_ROM_rdata_0 ) == ( 8'd46 )  ;
assign n2502____DOLLAR__6337 =  ( oc8051_ROM_rdata_0 ) == ( 8'd45 )  ;
assign n2503____DOLLAR__6341 =  ( oc8051_ROM_rdata_0 ) == ( 8'd44 )  ;
assign n2504____DOLLAR__6345 =  ( oc8051_ROM_rdata_0 ) == ( 8'd43 )  ;
assign n2505____DOLLAR__6349 =  ( oc8051_ROM_rdata_0 ) == ( 8'd42 )  ;
assign n2506____DOLLAR__6353 =  ( oc8051_ROM_rdata_0 ) == ( 8'd41 )  ;
assign n2507____DOLLAR__6357 =  ( oc8051_ROM_rdata_0 ) == ( 8'd40 )  ;
assign n2508____DOLLAR__6361 =  ( oc8051_ROM_rdata_0 ) == ( 8'd39 )  ;
assign n2509____DOLLAR__6365 =  ( oc8051_ROM_rdata_0 ) == ( 8'd38 )  ;
assign n2510____DOLLAR__6369 =  ( oc8051_ROM_rdata_0 ) == ( 8'd37 )  ;
assign n2511____DOLLAR__6373 =  ( oc8051_ROM_rdata_0 ) == ( 8'd36 )  ;
assign n2512____DOLLAR__6377 =  ( oc8051_ROM_rdata_0 ) == ( 8'd35 )  ;
assign n2513____DOLLAR__6381 =  ( oc8051_ROM_rdata_0 ) == ( 8'd34 )  ;
assign n2514____DOLLAR__6385 =  ( oc8051_ROM_rdata_0 ) == ( 8'd33 )  ;
assign n2515____DOLLAR__6389 =  ( oc8051_ROM_rdata_0 ) == ( 8'd32 )  ;
assign n2516____DOLLAR__6393 =  ( oc8051_ROM_rdata_0 ) == ( 8'd31 )  ;
assign n2517____DOLLAR__6397 =  ( oc8051_ROM_rdata_0 ) == ( 8'd30 )  ;
assign n2518____DOLLAR__6401 =  ( oc8051_ROM_rdata_0 ) == ( 8'd29 )  ;
assign n2519____DOLLAR__6405 =  ( oc8051_ROM_rdata_0 ) == ( 8'd28 )  ;
assign n2520____DOLLAR__6409 =  ( oc8051_ROM_rdata_0 ) == ( 8'd27 )  ;
assign n2521____DOLLAR__6413 =  ( oc8051_ROM_rdata_0 ) == ( 8'd26 )  ;
assign n2522____DOLLAR__6417 =  ( oc8051_ROM_rdata_0 ) == ( 8'd25 )  ;
assign n2523____DOLLAR__6421 =  ( oc8051_ROM_rdata_0 ) == ( 8'd24 )  ;
assign n2524____DOLLAR__6425 =  ( oc8051_ROM_rdata_0 ) == ( 8'd23 )  ;
assign n2525____DOLLAR__6429 =  ( oc8051_ROM_rdata_0 ) == ( 8'd22 )  ;
assign n2526____DOLLAR__6433 =  ( oc8051_ROM_rdata_0 ) == ( 8'd21 )  ;
assign n2527____DOLLAR__6437 =  ( oc8051_ROM_rdata_0 ) == ( 8'd20 )  ;
assign n2528____DOLLAR__6441 =  ( oc8051_ROM_rdata_0 ) == ( 8'd19 )  ;
assign n2529____DOLLAR__6445 =  ( oc8051_ROM_rdata_0 ) == ( 8'd18 )  ;
assign n2530____DOLLAR__6449 =  ( oc8051_ROM_rdata_0 ) == ( 8'd17 )  ;
assign n2531____DOLLAR__6453 =  ( oc8051_ROM_rdata_0 ) == ( 8'd16 )  ;
assign n2532____DOLLAR__6457 =  ( oc8051_ROM_rdata_0 ) == ( 8'd15 )  ;
assign n2533____DOLLAR__6461 =  ( oc8051_ROM_rdata_0 ) == ( 8'd14 )  ;
assign n2534____DOLLAR__6465 =  ( oc8051_ROM_rdata_0 ) == ( 8'd13 )  ;
assign n2535____DOLLAR__6469 =  ( oc8051_ROM_rdata_0 ) == ( 8'd12 )  ;
assign n2536____DOLLAR__6473 =  ( oc8051_ROM_rdata_0 ) == ( 8'd11 )  ;
assign n2537____DOLLAR__6477 =  ( oc8051_ROM_rdata_0 ) == ( 8'd10 )  ;
assign n2538____DOLLAR__6481 =  ( oc8051_ROM_rdata_0 ) == ( 8'd9 )  ;
assign n2539____DOLLAR__6485 =  ( oc8051_ROM_rdata_0 ) == ( 8'd8 )  ;
assign n2540____DOLLAR__6489 =  ( oc8051_ROM_rdata_0 ) == ( 8'd7 )  ;
assign n2541____DOLLAR__6493 =  ( oc8051_ROM_rdata_0 ) == ( 8'd6 )  ;
assign n2542____DOLLAR__6497 =  ( oc8051_ROM_rdata_0 ) == ( 8'd5 )  ;
assign n2543____DOLLAR__6501 =  ( oc8051_ROM_rdata_0 ) == ( 8'd4 )  ;
assign n2544____DOLLAR__6505 =  ( oc8051_ROM_rdata_0 ) == ( 8'd3 )  ;
assign n2545____DOLLAR__6509 =  ( oc8051_ROM_rdata_0 ) == ( 8'd2 )  ;
assign n2546____DOLLAR__6513 =  ( oc8051_ROM_rdata_0 ) == ( 8'd1 )  ;
assign n2547____DOLLAR__6517 =  ( oc8051_ROM_rdata_0 ) == ( 8'd0 )  ;
assign n2548____DOLLAR__6519 =  ( n2546____DOLLAR__6513 ) | ( n2547____DOLLAR__6517 )  ;
assign n2549____DOLLAR__6520 =  ( n2545____DOLLAR__6509 ) | ( n2548____DOLLAR__6519 )  ;
assign n2550____DOLLAR__6521 =  ( n2544____DOLLAR__6505 ) | ( n2549____DOLLAR__6520 )  ;
assign n2551____DOLLAR__6522 =  ( n2543____DOLLAR__6501 ) | ( n2550____DOLLAR__6521 )  ;
assign n2552____DOLLAR__6523 =  ( n2542____DOLLAR__6497 ) | ( n2551____DOLLAR__6522 )  ;
assign n2553____DOLLAR__6524 =  ( n2541____DOLLAR__6493 ) | ( n2552____DOLLAR__6523 )  ;
assign n2554____DOLLAR__6525 =  ( n2540____DOLLAR__6489 ) | ( n2553____DOLLAR__6524 )  ;
assign n2555____DOLLAR__6526 =  ( n2539____DOLLAR__6485 ) | ( n2554____DOLLAR__6525 )  ;
assign n2556____DOLLAR__6527 =  ( n2538____DOLLAR__6481 ) | ( n2555____DOLLAR__6526 )  ;
assign n2557____DOLLAR__6528 =  ( n2537____DOLLAR__6477 ) | ( n2556____DOLLAR__6527 )  ;
assign n2558____DOLLAR__6529 =  ( n2536____DOLLAR__6473 ) | ( n2557____DOLLAR__6528 )  ;
assign n2559____DOLLAR__6530 =  ( n2535____DOLLAR__6469 ) | ( n2558____DOLLAR__6529 )  ;
assign n2560____DOLLAR__6531 =  ( n2534____DOLLAR__6465 ) | ( n2559____DOLLAR__6530 )  ;
assign n2561____DOLLAR__6532 =  ( n2533____DOLLAR__6461 ) | ( n2560____DOLLAR__6531 )  ;
assign n2562____DOLLAR__6533 =  ( n2532____DOLLAR__6457 ) | ( n2561____DOLLAR__6532 )  ;
assign n2563____DOLLAR__6534 =  ( n2531____DOLLAR__6453 ) | ( n2562____DOLLAR__6533 )  ;
assign n2564____DOLLAR__6535 =  ( n2530____DOLLAR__6449 ) | ( n2563____DOLLAR__6534 )  ;
assign n2565____DOLLAR__6536 =  ( n2529____DOLLAR__6445 ) | ( n2564____DOLLAR__6535 )  ;
assign n2566____DOLLAR__6537 =  ( n2528____DOLLAR__6441 ) | ( n2565____DOLLAR__6536 )  ;
assign n2567____DOLLAR__6538 =  ( n2527____DOLLAR__6437 ) | ( n2566____DOLLAR__6537 )  ;
assign n2568____DOLLAR__6539 =  ( n2526____DOLLAR__6433 ) | ( n2567____DOLLAR__6538 )  ;
assign n2569____DOLLAR__6540 =  ( n2525____DOLLAR__6429 ) | ( n2568____DOLLAR__6539 )  ;
assign n2570____DOLLAR__6541 =  ( n2524____DOLLAR__6425 ) | ( n2569____DOLLAR__6540 )  ;
assign n2571____DOLLAR__6542 =  ( n2523____DOLLAR__6421 ) | ( n2570____DOLLAR__6541 )  ;
assign n2572____DOLLAR__6543 =  ( n2522____DOLLAR__6417 ) | ( n2571____DOLLAR__6542 )  ;
assign n2573____DOLLAR__6544 =  ( n2521____DOLLAR__6413 ) | ( n2572____DOLLAR__6543 )  ;
assign n2574____DOLLAR__6545 =  ( n2520____DOLLAR__6409 ) | ( n2573____DOLLAR__6544 )  ;
assign n2575____DOLLAR__6546 =  ( n2519____DOLLAR__6405 ) | ( n2574____DOLLAR__6545 )  ;
assign n2576____DOLLAR__6547 =  ( n2518____DOLLAR__6401 ) | ( n2575____DOLLAR__6546 )  ;
assign n2577____DOLLAR__6548 =  ( n2517____DOLLAR__6397 ) | ( n2576____DOLLAR__6547 )  ;
assign n2578____DOLLAR__6549 =  ( n2516____DOLLAR__6393 ) | ( n2577____DOLLAR__6548 )  ;
assign n2579____DOLLAR__6550 =  ( n2515____DOLLAR__6389 ) | ( n2578____DOLLAR__6549 )  ;
assign n2580____DOLLAR__6551 =  ( n2514____DOLLAR__6385 ) | ( n2579____DOLLAR__6550 )  ;
assign n2581____DOLLAR__6552 =  ( n2513____DOLLAR__6381 ) | ( n2580____DOLLAR__6551 )  ;
assign n2582____DOLLAR__6553 =  ( n2512____DOLLAR__6377 ) | ( n2581____DOLLAR__6552 )  ;
assign n2583____DOLLAR__6554 =  ( n2511____DOLLAR__6373 ) | ( n2582____DOLLAR__6553 )  ;
assign n2584____DOLLAR__6555 =  ( n2510____DOLLAR__6369 ) | ( n2583____DOLLAR__6554 )  ;
assign n2585____DOLLAR__6556 =  ( n2509____DOLLAR__6365 ) | ( n2584____DOLLAR__6555 )  ;
assign n2586____DOLLAR__6557 =  ( n2508____DOLLAR__6361 ) | ( n2585____DOLLAR__6556 )  ;
assign n2587____DOLLAR__6558 =  ( n2507____DOLLAR__6357 ) | ( n2586____DOLLAR__6557 )  ;
assign n2588____DOLLAR__6559 =  ( n2506____DOLLAR__6353 ) | ( n2587____DOLLAR__6558 )  ;
assign n2589____DOLLAR__6560 =  ( n2505____DOLLAR__6349 ) | ( n2588____DOLLAR__6559 )  ;
assign n2590____DOLLAR__6561 =  ( n2504____DOLLAR__6345 ) | ( n2589____DOLLAR__6560 )  ;
assign n2591____DOLLAR__6562 =  ( n2503____DOLLAR__6341 ) | ( n2590____DOLLAR__6561 )  ;
assign n2592____DOLLAR__6563 =  ( n2502____DOLLAR__6337 ) | ( n2591____DOLLAR__6562 )  ;
assign n2593____DOLLAR__6564 =  ( n2501____DOLLAR__6333 ) | ( n2592____DOLLAR__6563 )  ;
assign n2594____DOLLAR__6565 =  ( n2500____DOLLAR__6329 ) | ( n2593____DOLLAR__6564 )  ;
assign n2595____DOLLAR__6566 =  ( n2499____DOLLAR__6325 ) | ( n2594____DOLLAR__6565 )  ;
assign n2596____DOLLAR__6567 =  ( n2498____DOLLAR__6321 ) | ( n2595____DOLLAR__6566 )  ;
assign n2597____DOLLAR__6568 =  ( n2497____DOLLAR__6317 ) | ( n2596____DOLLAR__6567 )  ;
assign n2598____DOLLAR__6569 =  ( n2496____DOLLAR__6313 ) | ( n2597____DOLLAR__6568 )  ;
assign n2599____DOLLAR__6570 =  ( n2495____DOLLAR__6309 ) | ( n2598____DOLLAR__6569 )  ;
assign n2600____DOLLAR__6571 =  ( n2494____DOLLAR__6305 ) | ( n2599____DOLLAR__6570 )  ;
assign n2601____DOLLAR__6572 =  ( n2493____DOLLAR__6301 ) | ( n2600____DOLLAR__6571 )  ;
assign n2602____DOLLAR__6573 =  ( n2492____DOLLAR__6297 ) | ( n2601____DOLLAR__6572 )  ;
assign n2603____DOLLAR__6574 =  ( n2491____DOLLAR__6293 ) | ( n2602____DOLLAR__6573 )  ;
assign n2604____DOLLAR__6575 =  ( n2490____DOLLAR__6289 ) | ( n2603____DOLLAR__6574 )  ;
assign n2605____DOLLAR__6576 =  ( n2489____DOLLAR__6285 ) | ( n2604____DOLLAR__6575 )  ;
assign n2606____DOLLAR__6577 =  ( n2488____DOLLAR__6281 ) | ( n2605____DOLLAR__6576 )  ;
assign n2607____DOLLAR__6578 =  ( n2487____DOLLAR__6277 ) | ( n2606____DOLLAR__6577 )  ;
assign n2608____DOLLAR__6579 =  ( n2486____DOLLAR__6273 ) | ( n2607____DOLLAR__6578 )  ;
assign n2609____DOLLAR__6580 =  ( n2485____DOLLAR__6269 ) | ( n2608____DOLLAR__6579 )  ;
assign n2610____DOLLAR__6581 =  ( n2484____DOLLAR__6265 ) | ( n2609____DOLLAR__6580 )  ;
assign n2611____DOLLAR__6582 =  ( n2483____DOLLAR__6261 ) | ( n2610____DOLLAR__6581 )  ;
assign n2612____DOLLAR__6583 =  ( n2482____DOLLAR__6257 ) | ( n2611____DOLLAR__6582 )  ;
assign n2613____DOLLAR__6584 =  ( n2481____DOLLAR__6253 ) | ( n2612____DOLLAR__6583 )  ;
assign n2614____DOLLAR__6585 =  ( n2480____DOLLAR__6249 ) | ( n2613____DOLLAR__6584 )  ;
assign n2615____DOLLAR__6586 =  ( n2479____DOLLAR__6245 ) | ( n2614____DOLLAR__6585 )  ;
assign n2616____DOLLAR__6587 =  ( n2478____DOLLAR__6241 ) | ( n2615____DOLLAR__6586 )  ;
assign n2617____DOLLAR__6588 =  ( n2477____DOLLAR__6237 ) | ( n2616____DOLLAR__6587 )  ;
assign n2618____DOLLAR__6589 =  ( n2476____DOLLAR__6233 ) | ( n2617____DOLLAR__6588 )  ;
assign n2619____DOLLAR__6590 =  ( n2475____DOLLAR__6229 ) | ( n2618____DOLLAR__6589 )  ;
assign n2620____DOLLAR__6591 =  ( n2474____DOLLAR__6225 ) | ( n2619____DOLLAR__6590 )  ;
assign n2621____DOLLAR__6592 =  ( n2473____DOLLAR__6221 ) | ( n2620____DOLLAR__6591 )  ;
assign n2622____DOLLAR__6593 =  ( n2472____DOLLAR__6217 ) | ( n2621____DOLLAR__6592 )  ;
assign n2623____DOLLAR__6594 =  ( n2471____DOLLAR__6213 ) | ( n2622____DOLLAR__6593 )  ;
assign n2624____DOLLAR__6595 =  ( n2470____DOLLAR__6209 ) | ( n2623____DOLLAR__6594 )  ;
assign n2625____DOLLAR__6596 =  ( n2469____DOLLAR__6205 ) | ( n2624____DOLLAR__6595 )  ;
assign n2626____DOLLAR__6597 =  ( n2468____DOLLAR__6201 ) | ( n2625____DOLLAR__6596 )  ;
assign n2627____DOLLAR__6598 =  ( n2467____DOLLAR__6197 ) | ( n2626____DOLLAR__6597 )  ;
assign n2628____DOLLAR__6599 =  ( n2466____DOLLAR__6193 ) | ( n2627____DOLLAR__6598 )  ;
assign n2629____DOLLAR__6600 =  ( n2465____DOLLAR__6189 ) | ( n2628____DOLLAR__6599 )  ;
assign n2630____DOLLAR__6601 =  ( n2464____DOLLAR__6185 ) | ( n2629____DOLLAR__6600 )  ;
assign n2631____DOLLAR__6602 =  ( n2463____DOLLAR__6181 ) | ( n2630____DOLLAR__6601 )  ;
assign n2632____DOLLAR__6603 =  ( n2462____DOLLAR__6177 ) | ( n2631____DOLLAR__6602 )  ;
assign n2633____DOLLAR__6604 =  ( n2461____DOLLAR__6173 ) | ( n2632____DOLLAR__6603 )  ;
assign n2634____DOLLAR__6605 =  ( n2460____DOLLAR__6169 ) | ( n2633____DOLLAR__6604 )  ;
assign n2635____DOLLAR__6606 =  ( n2459____DOLLAR__6165 ) | ( n2634____DOLLAR__6605 )  ;
assign n2636____DOLLAR__6607 =  ( n2458____DOLLAR__6161 ) | ( n2635____DOLLAR__6606 )  ;
assign n2637____DOLLAR__6608 =  ( n2457____DOLLAR__6157 ) | ( n2636____DOLLAR__6607 )  ;
assign n2638____DOLLAR__6609 =  ( n2456____DOLLAR__6153 ) | ( n2637____DOLLAR__6608 )  ;
assign n2639____DOLLAR__6610 =  ( n2455____DOLLAR__6149 ) | ( n2638____DOLLAR__6609 )  ;
assign n2640____DOLLAR__6611 =  ( n2454____DOLLAR__6145 ) | ( n2639____DOLLAR__6610 )  ;
assign n2641____DOLLAR__6612 =  ( n2453____DOLLAR__6141 ) | ( n2640____DOLLAR__6611 )  ;
assign n2642____DOLLAR__6613 =  ( n2452____DOLLAR__6137 ) | ( n2641____DOLLAR__6612 )  ;
assign n2643____DOLLAR__6614 =  ( n2451____DOLLAR__6133 ) | ( n2642____DOLLAR__6613 )  ;
assign n2644____DOLLAR__6615 =  ( n2450____DOLLAR__6129 ) | ( n2643____DOLLAR__6614 )  ;
assign n2645____DOLLAR__6616 =  ( n2449____DOLLAR__6125 ) | ( n2644____DOLLAR__6615 )  ;
assign n2646____DOLLAR__6617 =  ( n2448____DOLLAR__6121 ) | ( n2645____DOLLAR__6616 )  ;
assign n2647____DOLLAR__6618 =  ( n2447____DOLLAR__6117 ) | ( n2646____DOLLAR__6617 )  ;
assign n2648____DOLLAR__6619 =  ( n2446____DOLLAR__6113 ) | ( n2647____DOLLAR__6618 )  ;
assign n2649____DOLLAR__6620 =  ( n2445____DOLLAR__6109 ) | ( n2648____DOLLAR__6619 )  ;
assign n2650____DOLLAR__6621 =  ( n2444____DOLLAR__6105 ) | ( n2649____DOLLAR__6620 )  ;
assign n2651____DOLLAR__6622 =  ( n2443____DOLLAR__6101 ) | ( n2650____DOLLAR__6621 )  ;
assign n2652____DOLLAR__6623 =  ( n2442____DOLLAR__6097 ) | ( n2651____DOLLAR__6622 )  ;
assign n2653____DOLLAR__6624 =  ( n2441____DOLLAR__6093 ) | ( n2652____DOLLAR__6623 )  ;
assign n2654____DOLLAR__6625 =  ( n2440____DOLLAR__6089 ) | ( n2653____DOLLAR__6624 )  ;
assign n2655____DOLLAR__6626 =  ( n2439____DOLLAR__6085 ) | ( n2654____DOLLAR__6625 )  ;
assign n2656____DOLLAR__6627 =  ( n2438____DOLLAR__6081 ) | ( n2655____DOLLAR__6626 )  ;
assign n2657____DOLLAR__6628 =  ( n2437____DOLLAR__6077 ) | ( n2656____DOLLAR__6627 )  ;
assign n2658____DOLLAR__6629 =  ( n2436____DOLLAR__6073 ) | ( n2657____DOLLAR__6628 )  ;
assign n2659____DOLLAR__6630 =  ( n2435____DOLLAR__6069 ) | ( n2658____DOLLAR__6629 )  ;
assign n2660____DOLLAR__6631 =  ( n2434____DOLLAR__6065 ) | ( n2659____DOLLAR__6630 )  ;
assign n2661____DOLLAR__6632 =  ( n2433____DOLLAR__6061 ) | ( n2660____DOLLAR__6631 )  ;
assign n2662____DOLLAR__6633 =  ( n2432____DOLLAR__6057 ) | ( n2661____DOLLAR__6632 )  ;
assign n2663____DOLLAR__6634 =  ( n2431____DOLLAR__6053 ) | ( n2662____DOLLAR__6633 )  ;
assign n2664____DOLLAR__6635 =  ( n2430____DOLLAR__6049 ) | ( n2663____DOLLAR__6634 )  ;
assign n2665____DOLLAR__6636 =  ( n2429____DOLLAR__6045 ) | ( n2664____DOLLAR__6635 )  ;
assign n2666____DOLLAR__6637 =  ( n2428____DOLLAR__6041 ) | ( n2665____DOLLAR__6636 )  ;
assign n2667____DOLLAR__6638 =  ( n2427____DOLLAR__6037 ) | ( n2666____DOLLAR__6637 )  ;
assign n2668____DOLLAR__6639 =  ( n2426____DOLLAR__6033 ) | ( n2667____DOLLAR__6638 )  ;
assign n2669____DOLLAR__6640 =  ( n2425____DOLLAR__6029 ) | ( n2668____DOLLAR__6639 )  ;
assign n2670____DOLLAR__6641 =  ( n2424____DOLLAR__6025 ) | ( n2669____DOLLAR__6640 )  ;
assign n2671____DOLLAR__6642 =  ( n2423____DOLLAR__6021 ) | ( n2670____DOLLAR__6641 )  ;
assign n2672____DOLLAR__6643 =  ( n2422____DOLLAR__6017 ) | ( n2671____DOLLAR__6642 )  ;
assign n2673____DOLLAR__6644 =  ( n2421____DOLLAR__6013 ) | ( n2672____DOLLAR__6643 )  ;
assign n2674____DOLLAR__6645 =  ( n2420____DOLLAR__6009 ) | ( n2673____DOLLAR__6644 )  ;
assign n2675____DOLLAR__6646 =  ( n2419____DOLLAR__6005 ) | ( n2674____DOLLAR__6645 )  ;
assign n2676____DOLLAR__6647 =  ( n2418____DOLLAR__6001 ) | ( n2675____DOLLAR__6646 )  ;
assign n2677____DOLLAR__6648 =  ( n2417____DOLLAR__5997 ) | ( n2676____DOLLAR__6647 )  ;
assign n2678____DOLLAR__6649 =  ( n2416____DOLLAR__5993 ) | ( n2677____DOLLAR__6648 )  ;
assign n2679____DOLLAR__6650 =  ( n2415____DOLLAR__5989 ) | ( n2678____DOLLAR__6649 )  ;
assign n2680____DOLLAR__6651 =  ( n2414____DOLLAR__5985 ) | ( n2679____DOLLAR__6650 )  ;
assign n2681____DOLLAR__6652 =  ( n2413____DOLLAR__5981 ) | ( n2680____DOLLAR__6651 )  ;
assign n2682____DOLLAR__6653 =  ( n2412____DOLLAR__5977 ) | ( n2681____DOLLAR__6652 )  ;
assign n2683____DOLLAR__6654 =  ( n2411____DOLLAR__5973 ) | ( n2682____DOLLAR__6653 )  ;
assign n2684____DOLLAR__6655 =  ( n2410____DOLLAR__5969 ) | ( n2683____DOLLAR__6654 )  ;
assign n2685____DOLLAR__6656 =  ( n2409____DOLLAR__5965 ) | ( n2684____DOLLAR__6655 )  ;
assign n2686____DOLLAR__6657 =  ( n2408____DOLLAR__5961 ) | ( n2685____DOLLAR__6656 )  ;
assign n2687____DOLLAR__6658 =  ( n2407____DOLLAR__5957 ) | ( n2686____DOLLAR__6657 )  ;
assign n2688____DOLLAR__6659 =  ( n2406____DOLLAR__5953 ) | ( n2687____DOLLAR__6658 )  ;
assign n2689____DOLLAR__6660 =  ( n2405____DOLLAR__5949 ) | ( n2688____DOLLAR__6659 )  ;
assign n2690____DOLLAR__6661 =  ( n2404____DOLLAR__5945 ) | ( n2689____DOLLAR__6660 )  ;
assign n2691____DOLLAR__6662 =  ( n2403____DOLLAR__5941 ) | ( n2690____DOLLAR__6661 )  ;
assign n2692____DOLLAR__6663 =  ( n2402____DOLLAR__5937 ) | ( n2691____DOLLAR__6662 )  ;
assign n2693____DOLLAR__6664 =  ( n2401____DOLLAR__5933 ) | ( n2692____DOLLAR__6663 )  ;
assign n2694____DOLLAR__6665 =  ( n2400____DOLLAR__5929 ) | ( n2693____DOLLAR__6664 )  ;
assign n2695____DOLLAR__6666 =  ( n2399____DOLLAR__5925 ) | ( n2694____DOLLAR__6665 )  ;
assign n2696____DOLLAR__6667 =  ( n2398____DOLLAR__5921 ) | ( n2695____DOLLAR__6666 )  ;
assign n2697____DOLLAR__6668 =  ( n2397____DOLLAR__5917 ) | ( n2696____DOLLAR__6667 )  ;
assign n2698____DOLLAR__6669 =  ( n2396____DOLLAR__5913 ) | ( n2697____DOLLAR__6668 )  ;
assign n2699____DOLLAR__6670 =  ( n2395____DOLLAR__5909 ) | ( n2698____DOLLAR__6669 )  ;
assign n2700____DOLLAR__6671 =  ( n2394____DOLLAR__5905 ) | ( n2699____DOLLAR__6670 )  ;
assign n2701____DOLLAR__6672 =  ( n2393____DOLLAR__5901 ) | ( n2700____DOLLAR__6671 )  ;
assign n2702____DOLLAR__6673 =  ( n2392____DOLLAR__5897 ) | ( n2701____DOLLAR__6672 )  ;
assign n2703____DOLLAR__6674 =  ( n2391____DOLLAR__5893 ) | ( n2702____DOLLAR__6673 )  ;
assign n2704____DOLLAR__6675 =  ( n2390____DOLLAR__5889 ) | ( n2703____DOLLAR__6674 )  ;
assign n2705____DOLLAR__6676 =  ( n2389____DOLLAR__5885 ) | ( n2704____DOLLAR__6675 )  ;
assign n2706____DOLLAR__6677 =  ( n2388____DOLLAR__5881 ) | ( n2705____DOLLAR__6676 )  ;
assign n2707____DOLLAR__6678 =  ( n2387____DOLLAR__5877 ) | ( n2706____DOLLAR__6677 )  ;
assign n2708____DOLLAR__6679 =  ( n2386____DOLLAR__5873 ) | ( n2707____DOLLAR__6678 )  ;
assign n2709____DOLLAR__6680 =  ( n2385____DOLLAR__5869 ) | ( n2708____DOLLAR__6679 )  ;
assign n2710____DOLLAR__6681 =  ( n2384____DOLLAR__5865 ) | ( n2709____DOLLAR__6680 )  ;
assign n2711____DOLLAR__6682 =  ( n2383____DOLLAR__5861 ) | ( n2710____DOLLAR__6681 )  ;
assign n2712____DOLLAR__6683 =  ( n2382____DOLLAR__5857 ) | ( n2711____DOLLAR__6682 )  ;
assign n2713____DOLLAR__6684 =  ( n2381____DOLLAR__5853 ) | ( n2712____DOLLAR__6683 )  ;
assign n2714____DOLLAR__6685 =  ( n2380____DOLLAR__5849 ) | ( n2713____DOLLAR__6684 )  ;
assign n2715____DOLLAR__6686 =  ( n2379____DOLLAR__5845 ) | ( n2714____DOLLAR__6685 )  ;
assign n2716____DOLLAR__6687 =  ( n2378____DOLLAR__5841 ) | ( n2715____DOLLAR__6686 )  ;
assign n2717____DOLLAR__6688 =  ( n2377____DOLLAR__5837 ) | ( n2716____DOLLAR__6687 )  ;
assign n2718____DOLLAR__6689 =  ( n2376____DOLLAR__5833 ) | ( n2717____DOLLAR__6688 )  ;
assign n2719____DOLLAR__6690 =  ( n2375____DOLLAR__5829 ) | ( n2718____DOLLAR__6689 )  ;
assign n2720____DOLLAR__6691 =  ( n2374____DOLLAR__5825 ) | ( n2719____DOLLAR__6690 )  ;
assign n2721____DOLLAR__6692 =  ( n2373____DOLLAR__5821 ) | ( n2720____DOLLAR__6691 )  ;
assign n2722____DOLLAR__6693 =  ( n2372____DOLLAR__5817 ) | ( n2721____DOLLAR__6692 )  ;
assign n2723____DOLLAR__6694 =  ( n2371____DOLLAR__5813 ) | ( n2722____DOLLAR__6693 )  ;
assign n2724____DOLLAR__6695 =  ( n2370____DOLLAR__5809 ) | ( n2723____DOLLAR__6694 )  ;
assign n2725____DOLLAR__6696 =  ( n2369____DOLLAR__5805 ) | ( n2724____DOLLAR__6695 )  ;
assign n2726____DOLLAR__6697 =  ( n2368____DOLLAR__5801 ) | ( n2725____DOLLAR__6696 )  ;
assign n2727____DOLLAR__6698 =  ( n2367____DOLLAR__5797 ) | ( n2726____DOLLAR__6697 )  ;
assign n2728____DOLLAR__6699 =  ( n2366____DOLLAR__5793 ) | ( n2727____DOLLAR__6698 )  ;
assign n2729____DOLLAR__6700 =  ( n2365____DOLLAR__5789 ) | ( n2728____DOLLAR__6699 )  ;
assign n2730____DOLLAR__6701 =  ( n2364____DOLLAR__5785 ) | ( n2729____DOLLAR__6700 )  ;
assign n2731____DOLLAR__6702 =  ( n2363____DOLLAR__5781 ) | ( n2730____DOLLAR__6701 )  ;
assign n2732____DOLLAR__6703 =  ( n2362____DOLLAR__5777 ) | ( n2731____DOLLAR__6702 )  ;
assign n2733____DOLLAR__6704 =  ( n2361____DOLLAR__5773 ) | ( n2732____DOLLAR__6703 )  ;
assign n2734____DOLLAR__6705 =  ( n2360____DOLLAR__5769 ) | ( n2733____DOLLAR__6704 )  ;
assign n2735____DOLLAR__6706 =  ( n2359____DOLLAR__5765 ) | ( n2734____DOLLAR__6705 )  ;
assign n2736____DOLLAR__6707 =  ( n2358____DOLLAR__5761 ) | ( n2735____DOLLAR__6706 )  ;
assign n2737____DOLLAR__6708 =  ( n2357____DOLLAR__5757 ) | ( n2736____DOLLAR__6707 )  ;
assign n2738____DOLLAR__6709 =  ( n2356____DOLLAR__5753 ) | ( n2737____DOLLAR__6708 )  ;
assign n2739____DOLLAR__6710 =  ( n2355____DOLLAR__5749 ) | ( n2738____DOLLAR__6709 )  ;
assign n2740____DOLLAR__6711 =  ( n2354____DOLLAR__5745 ) | ( n2739____DOLLAR__6710 )  ;
assign n2741____DOLLAR__6712 =  ( n2353____DOLLAR__5741 ) | ( n2740____DOLLAR__6711 )  ;
assign n2742____DOLLAR__6713 =  ( n2352____DOLLAR__5737 ) | ( n2741____DOLLAR__6712 )  ;
assign n2743____DOLLAR__6714 =  ( n2351____DOLLAR__5733 ) | ( n2742____DOLLAR__6713 )  ;
assign n2744____DOLLAR__6715 =  ( n2350____DOLLAR__5729 ) | ( n2743____DOLLAR__6714 )  ;
assign n2745____DOLLAR__6716 =  ( n2349____DOLLAR__5725 ) | ( n2744____DOLLAR__6715 )  ;
assign n2746____DOLLAR__6717 =  ( n2348____DOLLAR__5721 ) | ( n2745____DOLLAR__6716 )  ;
assign n2747____DOLLAR__6718 =  ( n2347____DOLLAR__5717 ) | ( n2746____DOLLAR__6717 )  ;
assign n2748____DOLLAR__6719 =  ( n2346____DOLLAR__5713 ) | ( n2747____DOLLAR__6718 )  ;
assign n2749____DOLLAR__6720 =  ( n2345____DOLLAR__5709 ) | ( n2748____DOLLAR__6719 )  ;
assign n2750____DOLLAR__6721 =  ( n2344____DOLLAR__5705 ) | ( n2749____DOLLAR__6720 )  ;
assign n2751____DOLLAR__6722 =  ( n2343____DOLLAR__5701 ) | ( n2750____DOLLAR__6721 )  ;
assign n2752____DOLLAR__6723 =  ( n2342____DOLLAR__5697 ) | ( n2751____DOLLAR__6722 )  ;
assign n2753____DOLLAR__6724 =  ( n2341____DOLLAR__5693 ) | ( n2752____DOLLAR__6723 )  ;
assign n2754____DOLLAR__6725 =  ( n2340____DOLLAR__5689 ) | ( n2753____DOLLAR__6724 )  ;
assign n2755____DOLLAR__6726 =  ( n2339____DOLLAR__5685 ) | ( n2754____DOLLAR__6725 )  ;
assign n2756____DOLLAR__6727 =  ( n2338____DOLLAR__5681 ) | ( n2755____DOLLAR__6726 )  ;
assign n2757____DOLLAR__6728 =  ( n2337____DOLLAR__5677 ) | ( n2756____DOLLAR__6727 )  ;
assign n2758____DOLLAR__6729 =  ( n2336____DOLLAR__5673 ) | ( n2757____DOLLAR__6728 )  ;
assign n2759____DOLLAR__6730 =  ( n2335____DOLLAR__5669 ) | ( n2758____DOLLAR__6729 )  ;
assign n2760____DOLLAR__6731 =  ( n2334____DOLLAR__5665 ) | ( n2759____DOLLAR__6730 )  ;
assign n2761____DOLLAR__6732 =  ( n2333____DOLLAR__5661 ) | ( n2760____DOLLAR__6731 )  ;
assign n2762____DOLLAR__6733 =  ( n2332____DOLLAR__5657 ) | ( n2761____DOLLAR__6732 )  ;
assign n2763____DOLLAR__6734 =  ( n2331____DOLLAR__5653 ) | ( n2762____DOLLAR__6733 )  ;
assign n2764____DOLLAR__6735 =  ( n2330____DOLLAR__5649 ) | ( n2763____DOLLAR__6734 )  ;
assign n2765____DOLLAR__6736 =  ( n2329____DOLLAR__5645 ) | ( n2764____DOLLAR__6735 )  ;
assign n2766____DOLLAR__6737 =  ( n2328____DOLLAR__5641 ) | ( n2765____DOLLAR__6736 )  ;
assign n2767____DOLLAR__6738 =  ( n2327____DOLLAR__5637 ) | ( n2766____DOLLAR__6737 )  ;
assign n2768____DOLLAR__6739 =  ( n2326____DOLLAR__5633 ) | ( n2767____DOLLAR__6738 )  ;
assign n2769____DOLLAR__6740 =  ( n2325____DOLLAR__5629 ) | ( n2768____DOLLAR__6739 )  ;
assign n2770____DOLLAR__6741 =  ( n2324____DOLLAR__5625 ) | ( n2769____DOLLAR__6740 )  ;
assign n2771____DOLLAR__6742 =  ( n2323____DOLLAR__5621 ) | ( n2770____DOLLAR__6741 )  ;
assign n2772____DOLLAR__6743 =  ( n2322____DOLLAR__5617 ) | ( n2771____DOLLAR__6742 )  ;
assign n2773____DOLLAR__6744 =  ( n2321____DOLLAR__5613 ) | ( n2772____DOLLAR__6743 )  ;
assign n2774____DOLLAR__6745 =  ( n2320____DOLLAR__5609 ) | ( n2773____DOLLAR__6744 )  ;
assign n2775____DOLLAR__6746 =  ( n2319____DOLLAR__5605 ) | ( n2774____DOLLAR__6745 )  ;
assign n2776____DOLLAR__6747 =  ( n2318____DOLLAR__5601 ) | ( n2775____DOLLAR__6746 )  ;
assign n2777____DOLLAR__6748 =  ( n2317____DOLLAR__5597 ) | ( n2776____DOLLAR__6747 )  ;
assign n2778____DOLLAR__6749 =  ( n2316____DOLLAR__5593 ) | ( n2777____DOLLAR__6748 )  ;
assign n2779____DOLLAR__6750 =  ( n2315____DOLLAR__5589 ) | ( n2778____DOLLAR__6749 )  ;
assign n2780____DOLLAR__6751 =  ( n2314____DOLLAR__5585 ) | ( n2779____DOLLAR__6750 )  ;
assign n2781____DOLLAR__6752 =  ( n2313____DOLLAR__5581 ) | ( n2780____DOLLAR__6751 )  ;
assign n2782____DOLLAR__6753 =  ( n2312____DOLLAR__5577 ) | ( n2781____DOLLAR__6752 )  ;
assign n2783____DOLLAR__6754 =  ( n2311____DOLLAR__5573 ) | ( n2782____DOLLAR__6753 )  ;
assign n2784____DOLLAR__6755 =  ( n2310____DOLLAR__5569 ) | ( n2783____DOLLAR__6754 )  ;
assign n2785____DOLLAR__6756 =  ( n2309____DOLLAR__5565 ) | ( n2784____DOLLAR__6755 )  ;
assign n2786____DOLLAR__6757 =  ( n2308____DOLLAR__5561 ) | ( n2785____DOLLAR__6756 )  ;
assign n2787____DOLLAR__6758 =  ( n2307____DOLLAR__5557 ) | ( n2786____DOLLAR__6757 )  ;
assign n2788____DOLLAR__6759 =  ( n2306____DOLLAR__5553 ) | ( n2787____DOLLAR__6758 )  ;
assign n2789____DOLLAR__6760 =  ( n2305____DOLLAR__5549 ) | ( n2788____DOLLAR__6759 )  ;
assign n2790____DOLLAR__6761 =  ( n2304____DOLLAR__5545 ) | ( n2789____DOLLAR__6760 )  ;
assign n2791____DOLLAR__6762 =  ( n2303____DOLLAR__5541 ) | ( n2790____DOLLAR__6761 )  ;
assign n2792____DOLLAR__6763 =  ( n2302____DOLLAR__5537 ) | ( n2791____DOLLAR__6762 )  ;
assign n2793____DOLLAR__6764 =  ( n2301____DOLLAR__5533 ) | ( n2792____DOLLAR__6763 )  ;
assign n2794____DOLLAR__6765 =  ( n2300____DOLLAR__5529 ) | ( n2793____DOLLAR__6764 )  ;
assign n2795____DOLLAR__6766 =  ( n2299____DOLLAR__5525 ) | ( n2794____DOLLAR__6765 )  ;
assign n2796____DOLLAR__6767 =  ( n2298____DOLLAR__5521 ) | ( n2795____DOLLAR__6766 )  ;
assign n2797____DOLLAR__6770 =  ( n2796____DOLLAR__6767 ) ? ( 16'd0 ) : ( XRAM_ADDR ) ;
assign n2798____DOLLAR__6771 =  ( n2296____DOLLAR__5510 ) ? ( n2297____DOLLAR__5515 ) : ( n2797____DOLLAR__6770 ) ;
assign n2799____DOLLAR__6772 =  ( n2256____DOLLAR__5471 ) ? ( n2293____DOLLAR__5498 ) : ( n2798____DOLLAR__6771 ) ;
assign n2800____DOLLAR__6773 =  ( n2216____DOLLAR__5432 ) ? ( n2253____DOLLAR__5459 ) : ( n2799____DOLLAR__6772 ) ;
assign n2801____DOLLAR__6778 =  ( oc8051_ROM_rdata_0 ) == ( 8'd243 )  ;
assign n2802____DOLLAR__6782 =  ( oc8051_ROM_rdata_0 ) == ( 8'd242 )  ;
assign n2803____DOLLAR__6786 =  ( oc8051_ROM_rdata_0 ) == ( 8'd240 )  ;
assign n2804____DOLLAR__6788 =  ( n2802____DOLLAR__6782 ) | ( n2803____DOLLAR__6786 )  ;
assign n2805____DOLLAR__6789 =  ( n2801____DOLLAR__6778 ) | ( n2804____DOLLAR__6788 )  ;
assign n2806____DOLLAR__6794 =  ( oc8051_ROM_rdata_0 ) == ( 8'd255 )  ;
assign n2807____DOLLAR__6798 =  ( oc8051_ROM_rdata_0 ) == ( 8'd254 )  ;
assign n2808____DOLLAR__6802 =  ( oc8051_ROM_rdata_0 ) == ( 8'd253 )  ;
assign n2809____DOLLAR__6806 =  ( oc8051_ROM_rdata_0 ) == ( 8'd252 )  ;
assign n2810____DOLLAR__6810 =  ( oc8051_ROM_rdata_0 ) == ( 8'd251 )  ;
assign n2811____DOLLAR__6814 =  ( oc8051_ROM_rdata_0 ) == ( 8'd250 )  ;
assign n2812____DOLLAR__6818 =  ( oc8051_ROM_rdata_0 ) == ( 8'd249 )  ;
assign n2813____DOLLAR__6822 =  ( oc8051_ROM_rdata_0 ) == ( 8'd248 )  ;
assign n2814____DOLLAR__6826 =  ( oc8051_ROM_rdata_0 ) == ( 8'd247 )  ;
assign n2815____DOLLAR__6830 =  ( oc8051_ROM_rdata_0 ) == ( 8'd246 )  ;
assign n2816____DOLLAR__6834 =  ( oc8051_ROM_rdata_0 ) == ( 8'd245 )  ;
assign n2817____DOLLAR__6838 =  ( oc8051_ROM_rdata_0 ) == ( 8'd244 )  ;
assign n2818____DOLLAR__6842 =  ( oc8051_ROM_rdata_0 ) == ( 8'd241 )  ;
assign n2819____DOLLAR__6846 =  ( oc8051_ROM_rdata_0 ) == ( 8'd239 )  ;
assign n2820____DOLLAR__6850 =  ( oc8051_ROM_rdata_0 ) == ( 8'd238 )  ;
assign n2821____DOLLAR__6854 =  ( oc8051_ROM_rdata_0 ) == ( 8'd237 )  ;
assign n2822____DOLLAR__6858 =  ( oc8051_ROM_rdata_0 ) == ( 8'd236 )  ;
assign n2823____DOLLAR__6862 =  ( oc8051_ROM_rdata_0 ) == ( 8'd235 )  ;
assign n2824____DOLLAR__6866 =  ( oc8051_ROM_rdata_0 ) == ( 8'd234 )  ;
assign n2825____DOLLAR__6870 =  ( oc8051_ROM_rdata_0 ) == ( 8'd233 )  ;
assign n2826____DOLLAR__6874 =  ( oc8051_ROM_rdata_0 ) == ( 8'd232 )  ;
assign n2827____DOLLAR__6878 =  ( oc8051_ROM_rdata_0 ) == ( 8'd231 )  ;
assign n2828____DOLLAR__6882 =  ( oc8051_ROM_rdata_0 ) == ( 8'd230 )  ;
assign n2829____DOLLAR__6886 =  ( oc8051_ROM_rdata_0 ) == ( 8'd229 )  ;
assign n2830____DOLLAR__6890 =  ( oc8051_ROM_rdata_0 ) == ( 8'd228 )  ;
assign n2831____DOLLAR__6894 =  ( oc8051_ROM_rdata_0 ) == ( 8'd227 )  ;
assign n2832____DOLLAR__6898 =  ( oc8051_ROM_rdata_0 ) == ( 8'd226 )  ;
assign n2833____DOLLAR__6902 =  ( oc8051_ROM_rdata_0 ) == ( 8'd225 )  ;
assign n2834____DOLLAR__6906 =  ( oc8051_ROM_rdata_0 ) == ( 8'd224 )  ;
assign n2835____DOLLAR__6910 =  ( oc8051_ROM_rdata_0 ) == ( 8'd223 )  ;
assign n2836____DOLLAR__6914 =  ( oc8051_ROM_rdata_0 ) == ( 8'd222 )  ;
assign n2837____DOLLAR__6918 =  ( oc8051_ROM_rdata_0 ) == ( 8'd221 )  ;
assign n2838____DOLLAR__6922 =  ( oc8051_ROM_rdata_0 ) == ( 8'd220 )  ;
assign n2839____DOLLAR__6926 =  ( oc8051_ROM_rdata_0 ) == ( 8'd219 )  ;
assign n2840____DOLLAR__6930 =  ( oc8051_ROM_rdata_0 ) == ( 8'd218 )  ;
assign n2841____DOLLAR__6934 =  ( oc8051_ROM_rdata_0 ) == ( 8'd217 )  ;
assign n2842____DOLLAR__6938 =  ( oc8051_ROM_rdata_0 ) == ( 8'd216 )  ;
assign n2843____DOLLAR__6942 =  ( oc8051_ROM_rdata_0 ) == ( 8'd215 )  ;
assign n2844____DOLLAR__6946 =  ( oc8051_ROM_rdata_0 ) == ( 8'd214 )  ;
assign n2845____DOLLAR__6950 =  ( oc8051_ROM_rdata_0 ) == ( 8'd213 )  ;
assign n2846____DOLLAR__6954 =  ( oc8051_ROM_rdata_0 ) == ( 8'd212 )  ;
assign n2847____DOLLAR__6958 =  ( oc8051_ROM_rdata_0 ) == ( 8'd211 )  ;
assign n2848____DOLLAR__6962 =  ( oc8051_ROM_rdata_0 ) == ( 8'd210 )  ;
assign n2849____DOLLAR__6966 =  ( oc8051_ROM_rdata_0 ) == ( 8'd209 )  ;
assign n2850____DOLLAR__6970 =  ( oc8051_ROM_rdata_0 ) == ( 8'd208 )  ;
assign n2851____DOLLAR__6974 =  ( oc8051_ROM_rdata_0 ) == ( 8'd207 )  ;
assign n2852____DOLLAR__6978 =  ( oc8051_ROM_rdata_0 ) == ( 8'd206 )  ;
assign n2853____DOLLAR__6982 =  ( oc8051_ROM_rdata_0 ) == ( 8'd205 )  ;
assign n2854____DOLLAR__6986 =  ( oc8051_ROM_rdata_0 ) == ( 8'd204 )  ;
assign n2855____DOLLAR__6990 =  ( oc8051_ROM_rdata_0 ) == ( 8'd203 )  ;
assign n2856____DOLLAR__6994 =  ( oc8051_ROM_rdata_0 ) == ( 8'd202 )  ;
assign n2857____DOLLAR__6998 =  ( oc8051_ROM_rdata_0 ) == ( 8'd201 )  ;
assign n2858____DOLLAR__7002 =  ( oc8051_ROM_rdata_0 ) == ( 8'd200 )  ;
assign n2859____DOLLAR__7006 =  ( oc8051_ROM_rdata_0 ) == ( 8'd199 )  ;
assign n2860____DOLLAR__7010 =  ( oc8051_ROM_rdata_0 ) == ( 8'd198 )  ;
assign n2861____DOLLAR__7014 =  ( oc8051_ROM_rdata_0 ) == ( 8'd197 )  ;
assign n2862____DOLLAR__7018 =  ( oc8051_ROM_rdata_0 ) == ( 8'd196 )  ;
assign n2863____DOLLAR__7022 =  ( oc8051_ROM_rdata_0 ) == ( 8'd195 )  ;
assign n2864____DOLLAR__7026 =  ( oc8051_ROM_rdata_0 ) == ( 8'd194 )  ;
assign n2865____DOLLAR__7030 =  ( oc8051_ROM_rdata_0 ) == ( 8'd193 )  ;
assign n2866____DOLLAR__7034 =  ( oc8051_ROM_rdata_0 ) == ( 8'd192 )  ;
assign n2867____DOLLAR__7038 =  ( oc8051_ROM_rdata_0 ) == ( 8'd191 )  ;
assign n2868____DOLLAR__7042 =  ( oc8051_ROM_rdata_0 ) == ( 8'd190 )  ;
assign n2869____DOLLAR__7046 =  ( oc8051_ROM_rdata_0 ) == ( 8'd189 )  ;
assign n2870____DOLLAR__7050 =  ( oc8051_ROM_rdata_0 ) == ( 8'd188 )  ;
assign n2871____DOLLAR__7054 =  ( oc8051_ROM_rdata_0 ) == ( 8'd187 )  ;
assign n2872____DOLLAR__7058 =  ( oc8051_ROM_rdata_0 ) == ( 8'd186 )  ;
assign n2873____DOLLAR__7062 =  ( oc8051_ROM_rdata_0 ) == ( 8'd185 )  ;
assign n2874____DOLLAR__7066 =  ( oc8051_ROM_rdata_0 ) == ( 8'd184 )  ;
assign n2875____DOLLAR__7070 =  ( oc8051_ROM_rdata_0 ) == ( 8'd183 )  ;
assign n2876____DOLLAR__7074 =  ( oc8051_ROM_rdata_0 ) == ( 8'd182 )  ;
assign n2877____DOLLAR__7078 =  ( oc8051_ROM_rdata_0 ) == ( 8'd181 )  ;
assign n2878____DOLLAR__7082 =  ( oc8051_ROM_rdata_0 ) == ( 8'd180 )  ;
assign n2879____DOLLAR__7086 =  ( oc8051_ROM_rdata_0 ) == ( 8'd179 )  ;
assign n2880____DOLLAR__7090 =  ( oc8051_ROM_rdata_0 ) == ( 8'd178 )  ;
assign n2881____DOLLAR__7094 =  ( oc8051_ROM_rdata_0 ) == ( 8'd177 )  ;
assign n2882____DOLLAR__7098 =  ( oc8051_ROM_rdata_0 ) == ( 8'd176 )  ;
assign n2883____DOLLAR__7102 =  ( oc8051_ROM_rdata_0 ) == ( 8'd175 )  ;
assign n2884____DOLLAR__7106 =  ( oc8051_ROM_rdata_0 ) == ( 8'd174 )  ;
assign n2885____DOLLAR__7110 =  ( oc8051_ROM_rdata_0 ) == ( 8'd173 )  ;
assign n2886____DOLLAR__7114 =  ( oc8051_ROM_rdata_0 ) == ( 8'd172 )  ;
assign n2887____DOLLAR__7118 =  ( oc8051_ROM_rdata_0 ) == ( 8'd171 )  ;
assign n2888____DOLLAR__7122 =  ( oc8051_ROM_rdata_0 ) == ( 8'd170 )  ;
assign n2889____DOLLAR__7126 =  ( oc8051_ROM_rdata_0 ) == ( 8'd169 )  ;
assign n2890____DOLLAR__7130 =  ( oc8051_ROM_rdata_0 ) == ( 8'd168 )  ;
assign n2891____DOLLAR__7134 =  ( oc8051_ROM_rdata_0 ) == ( 8'd167 )  ;
assign n2892____DOLLAR__7138 =  ( oc8051_ROM_rdata_0 ) == ( 8'd166 )  ;
assign n2893____DOLLAR__7142 =  ( oc8051_ROM_rdata_0 ) == ( 8'd165 )  ;
assign n2894____DOLLAR__7146 =  ( oc8051_ROM_rdata_0 ) == ( 8'd164 )  ;
assign n2895____DOLLAR__7150 =  ( oc8051_ROM_rdata_0 ) == ( 8'd163 )  ;
assign n2896____DOLLAR__7154 =  ( oc8051_ROM_rdata_0 ) == ( 8'd162 )  ;
assign n2897____DOLLAR__7158 =  ( oc8051_ROM_rdata_0 ) == ( 8'd161 )  ;
assign n2898____DOLLAR__7162 =  ( oc8051_ROM_rdata_0 ) == ( 8'd160 )  ;
assign n2899____DOLLAR__7166 =  ( oc8051_ROM_rdata_0 ) == ( 8'd159 )  ;
assign n2900____DOLLAR__7170 =  ( oc8051_ROM_rdata_0 ) == ( 8'd158 )  ;
assign n2901____DOLLAR__7174 =  ( oc8051_ROM_rdata_0 ) == ( 8'd157 )  ;
assign n2902____DOLLAR__7178 =  ( oc8051_ROM_rdata_0 ) == ( 8'd156 )  ;
assign n2903____DOLLAR__7182 =  ( oc8051_ROM_rdata_0 ) == ( 8'd155 )  ;
assign n2904____DOLLAR__7186 =  ( oc8051_ROM_rdata_0 ) == ( 8'd154 )  ;
assign n2905____DOLLAR__7190 =  ( oc8051_ROM_rdata_0 ) == ( 8'd153 )  ;
assign n2906____DOLLAR__7194 =  ( oc8051_ROM_rdata_0 ) == ( 8'd152 )  ;
assign n2907____DOLLAR__7198 =  ( oc8051_ROM_rdata_0 ) == ( 8'd151 )  ;
assign n2908____DOLLAR__7202 =  ( oc8051_ROM_rdata_0 ) == ( 8'd150 )  ;
assign n2909____DOLLAR__7206 =  ( oc8051_ROM_rdata_0 ) == ( 8'd149 )  ;
assign n2910____DOLLAR__7210 =  ( oc8051_ROM_rdata_0 ) == ( 8'd148 )  ;
assign n2911____DOLLAR__7214 =  ( oc8051_ROM_rdata_0 ) == ( 8'd147 )  ;
assign n2912____DOLLAR__7218 =  ( oc8051_ROM_rdata_0 ) == ( 8'd146 )  ;
assign n2913____DOLLAR__7222 =  ( oc8051_ROM_rdata_0 ) == ( 8'd145 )  ;
assign n2914____DOLLAR__7226 =  ( oc8051_ROM_rdata_0 ) == ( 8'd144 )  ;
assign n2915____DOLLAR__7230 =  ( oc8051_ROM_rdata_0 ) == ( 8'd143 )  ;
assign n2916____DOLLAR__7234 =  ( oc8051_ROM_rdata_0 ) == ( 8'd142 )  ;
assign n2917____DOLLAR__7238 =  ( oc8051_ROM_rdata_0 ) == ( 8'd141 )  ;
assign n2918____DOLLAR__7242 =  ( oc8051_ROM_rdata_0 ) == ( 8'd140 )  ;
assign n2919____DOLLAR__7246 =  ( oc8051_ROM_rdata_0 ) == ( 8'd139 )  ;
assign n2920____DOLLAR__7250 =  ( oc8051_ROM_rdata_0 ) == ( 8'd138 )  ;
assign n2921____DOLLAR__7254 =  ( oc8051_ROM_rdata_0 ) == ( 8'd137 )  ;
assign n2922____DOLLAR__7258 =  ( oc8051_ROM_rdata_0 ) == ( 8'd136 )  ;
assign n2923____DOLLAR__7262 =  ( oc8051_ROM_rdata_0 ) == ( 8'd135 )  ;
assign n2924____DOLLAR__7266 =  ( oc8051_ROM_rdata_0 ) == ( 8'd134 )  ;
assign n2925____DOLLAR__7270 =  ( oc8051_ROM_rdata_0 ) == ( 8'd133 )  ;
assign n2926____DOLLAR__7274 =  ( oc8051_ROM_rdata_0 ) == ( 8'd132 )  ;
assign n2927____DOLLAR__7278 =  ( oc8051_ROM_rdata_0 ) == ( 8'd131 )  ;
assign n2928____DOLLAR__7282 =  ( oc8051_ROM_rdata_0 ) == ( 8'd130 )  ;
assign n2929____DOLLAR__7286 =  ( oc8051_ROM_rdata_0 ) == ( 8'd129 )  ;
assign n2930____DOLLAR__7290 =  ( oc8051_ROM_rdata_0 ) == ( 8'd128 )  ;
assign n2931____DOLLAR__7294 =  ( oc8051_ROM_rdata_0 ) == ( 8'd127 )  ;
assign n2932____DOLLAR__7298 =  ( oc8051_ROM_rdata_0 ) == ( 8'd126 )  ;
assign n2933____DOLLAR__7302 =  ( oc8051_ROM_rdata_0 ) == ( 8'd125 )  ;
assign n2934____DOLLAR__7306 =  ( oc8051_ROM_rdata_0 ) == ( 8'd124 )  ;
assign n2935____DOLLAR__7310 =  ( oc8051_ROM_rdata_0 ) == ( 8'd123 )  ;
assign n2936____DOLLAR__7314 =  ( oc8051_ROM_rdata_0 ) == ( 8'd122 )  ;
assign n2937____DOLLAR__7318 =  ( oc8051_ROM_rdata_0 ) == ( 8'd121 )  ;
assign n2938____DOLLAR__7322 =  ( oc8051_ROM_rdata_0 ) == ( 8'd120 )  ;
assign n2939____DOLLAR__7326 =  ( oc8051_ROM_rdata_0 ) == ( 8'd119 )  ;
assign n2940____DOLLAR__7330 =  ( oc8051_ROM_rdata_0 ) == ( 8'd118 )  ;
assign n2941____DOLLAR__7334 =  ( oc8051_ROM_rdata_0 ) == ( 8'd117 )  ;
assign n2942____DOLLAR__7338 =  ( oc8051_ROM_rdata_0 ) == ( 8'd116 )  ;
assign n2943____DOLLAR__7342 =  ( oc8051_ROM_rdata_0 ) == ( 8'd115 )  ;
assign n2944____DOLLAR__7346 =  ( oc8051_ROM_rdata_0 ) == ( 8'd114 )  ;
assign n2945____DOLLAR__7350 =  ( oc8051_ROM_rdata_0 ) == ( 8'd113 )  ;
assign n2946____DOLLAR__7354 =  ( oc8051_ROM_rdata_0 ) == ( 8'd112 )  ;
assign n2947____DOLLAR__7358 =  ( oc8051_ROM_rdata_0 ) == ( 8'd111 )  ;
assign n2948____DOLLAR__7362 =  ( oc8051_ROM_rdata_0 ) == ( 8'd110 )  ;
assign n2949____DOLLAR__7366 =  ( oc8051_ROM_rdata_0 ) == ( 8'd109 )  ;
assign n2950____DOLLAR__7370 =  ( oc8051_ROM_rdata_0 ) == ( 8'd108 )  ;
assign n2951____DOLLAR__7374 =  ( oc8051_ROM_rdata_0 ) == ( 8'd107 )  ;
assign n2952____DOLLAR__7378 =  ( oc8051_ROM_rdata_0 ) == ( 8'd106 )  ;
assign n2953____DOLLAR__7382 =  ( oc8051_ROM_rdata_0 ) == ( 8'd105 )  ;
assign n2954____DOLLAR__7386 =  ( oc8051_ROM_rdata_0 ) == ( 8'd104 )  ;
assign n2955____DOLLAR__7390 =  ( oc8051_ROM_rdata_0 ) == ( 8'd103 )  ;
assign n2956____DOLLAR__7394 =  ( oc8051_ROM_rdata_0 ) == ( 8'd102 )  ;
assign n2957____DOLLAR__7398 =  ( oc8051_ROM_rdata_0 ) == ( 8'd101 )  ;
assign n2958____DOLLAR__7402 =  ( oc8051_ROM_rdata_0 ) == ( 8'd100 )  ;
assign n2959____DOLLAR__7406 =  ( oc8051_ROM_rdata_0 ) == ( 8'd99 )  ;
assign n2960____DOLLAR__7410 =  ( oc8051_ROM_rdata_0 ) == ( 8'd98 )  ;
assign n2961____DOLLAR__7414 =  ( oc8051_ROM_rdata_0 ) == ( 8'd97 )  ;
assign n2962____DOLLAR__7418 =  ( oc8051_ROM_rdata_0 ) == ( 8'd96 )  ;
assign n2963____DOLLAR__7422 =  ( oc8051_ROM_rdata_0 ) == ( 8'd95 )  ;
assign n2964____DOLLAR__7426 =  ( oc8051_ROM_rdata_0 ) == ( 8'd94 )  ;
assign n2965____DOLLAR__7430 =  ( oc8051_ROM_rdata_0 ) == ( 8'd93 )  ;
assign n2966____DOLLAR__7434 =  ( oc8051_ROM_rdata_0 ) == ( 8'd92 )  ;
assign n2967____DOLLAR__7438 =  ( oc8051_ROM_rdata_0 ) == ( 8'd91 )  ;
assign n2968____DOLLAR__7442 =  ( oc8051_ROM_rdata_0 ) == ( 8'd90 )  ;
assign n2969____DOLLAR__7446 =  ( oc8051_ROM_rdata_0 ) == ( 8'd89 )  ;
assign n2970____DOLLAR__7450 =  ( oc8051_ROM_rdata_0 ) == ( 8'd88 )  ;
assign n2971____DOLLAR__7454 =  ( oc8051_ROM_rdata_0 ) == ( 8'd87 )  ;
assign n2972____DOLLAR__7458 =  ( oc8051_ROM_rdata_0 ) == ( 8'd86 )  ;
assign n2973____DOLLAR__7462 =  ( oc8051_ROM_rdata_0 ) == ( 8'd85 )  ;
assign n2974____DOLLAR__7466 =  ( oc8051_ROM_rdata_0 ) == ( 8'd84 )  ;
assign n2975____DOLLAR__7470 =  ( oc8051_ROM_rdata_0 ) == ( 8'd83 )  ;
assign n2976____DOLLAR__7474 =  ( oc8051_ROM_rdata_0 ) == ( 8'd82 )  ;
assign n2977____DOLLAR__7478 =  ( oc8051_ROM_rdata_0 ) == ( 8'd81 )  ;
assign n2978____DOLLAR__7482 =  ( oc8051_ROM_rdata_0 ) == ( 8'd80 )  ;
assign n2979____DOLLAR__7486 =  ( oc8051_ROM_rdata_0 ) == ( 8'd79 )  ;
assign n2980____DOLLAR__7490 =  ( oc8051_ROM_rdata_0 ) == ( 8'd78 )  ;
assign n2981____DOLLAR__7494 =  ( oc8051_ROM_rdata_0 ) == ( 8'd77 )  ;
assign n2982____DOLLAR__7498 =  ( oc8051_ROM_rdata_0 ) == ( 8'd76 )  ;
assign n2983____DOLLAR__7502 =  ( oc8051_ROM_rdata_0 ) == ( 8'd75 )  ;
assign n2984____DOLLAR__7506 =  ( oc8051_ROM_rdata_0 ) == ( 8'd74 )  ;
assign n2985____DOLLAR__7510 =  ( oc8051_ROM_rdata_0 ) == ( 8'd73 )  ;
assign n2986____DOLLAR__7514 =  ( oc8051_ROM_rdata_0 ) == ( 8'd72 )  ;
assign n2987____DOLLAR__7518 =  ( oc8051_ROM_rdata_0 ) == ( 8'd71 )  ;
assign n2988____DOLLAR__7522 =  ( oc8051_ROM_rdata_0 ) == ( 8'd70 )  ;
assign n2989____DOLLAR__7526 =  ( oc8051_ROM_rdata_0 ) == ( 8'd69 )  ;
assign n2990____DOLLAR__7530 =  ( oc8051_ROM_rdata_0 ) == ( 8'd68 )  ;
assign n2991____DOLLAR__7534 =  ( oc8051_ROM_rdata_0 ) == ( 8'd67 )  ;
assign n2992____DOLLAR__7538 =  ( oc8051_ROM_rdata_0 ) == ( 8'd66 )  ;
assign n2993____DOLLAR__7542 =  ( oc8051_ROM_rdata_0 ) == ( 8'd65 )  ;
assign n2994____DOLLAR__7546 =  ( oc8051_ROM_rdata_0 ) == ( 8'd64 )  ;
assign n2995____DOLLAR__7550 =  ( oc8051_ROM_rdata_0 ) == ( 8'd63 )  ;
assign n2996____DOLLAR__7554 =  ( oc8051_ROM_rdata_0 ) == ( 8'd62 )  ;
assign n2997____DOLLAR__7558 =  ( oc8051_ROM_rdata_0 ) == ( 8'd61 )  ;
assign n2998____DOLLAR__7562 =  ( oc8051_ROM_rdata_0 ) == ( 8'd60 )  ;
assign n2999____DOLLAR__7566 =  ( oc8051_ROM_rdata_0 ) == ( 8'd59 )  ;
assign n3000____DOLLAR__7570 =  ( oc8051_ROM_rdata_0 ) == ( 8'd58 )  ;
assign n3001____DOLLAR__7574 =  ( oc8051_ROM_rdata_0 ) == ( 8'd57 )  ;
assign n3002____DOLLAR__7578 =  ( oc8051_ROM_rdata_0 ) == ( 8'd56 )  ;
assign n3003____DOLLAR__7582 =  ( oc8051_ROM_rdata_0 ) == ( 8'd55 )  ;
assign n3004____DOLLAR__7586 =  ( oc8051_ROM_rdata_0 ) == ( 8'd54 )  ;
assign n3005____DOLLAR__7590 =  ( oc8051_ROM_rdata_0 ) == ( 8'd53 )  ;
assign n3006____DOLLAR__7594 =  ( oc8051_ROM_rdata_0 ) == ( 8'd52 )  ;
assign n3007____DOLLAR__7598 =  ( oc8051_ROM_rdata_0 ) == ( 8'd51 )  ;
assign n3008____DOLLAR__7602 =  ( oc8051_ROM_rdata_0 ) == ( 8'd50 )  ;
assign n3009____DOLLAR__7606 =  ( oc8051_ROM_rdata_0 ) == ( 8'd49 )  ;
assign n3010____DOLLAR__7610 =  ( oc8051_ROM_rdata_0 ) == ( 8'd48 )  ;
assign n3011____DOLLAR__7614 =  ( oc8051_ROM_rdata_0 ) == ( 8'd47 )  ;
assign n3012____DOLLAR__7618 =  ( oc8051_ROM_rdata_0 ) == ( 8'd46 )  ;
assign n3013____DOLLAR__7622 =  ( oc8051_ROM_rdata_0 ) == ( 8'd45 )  ;
assign n3014____DOLLAR__7626 =  ( oc8051_ROM_rdata_0 ) == ( 8'd44 )  ;
assign n3015____DOLLAR__7630 =  ( oc8051_ROM_rdata_0 ) == ( 8'd43 )  ;
assign n3016____DOLLAR__7634 =  ( oc8051_ROM_rdata_0 ) == ( 8'd42 )  ;
assign n3017____DOLLAR__7638 =  ( oc8051_ROM_rdata_0 ) == ( 8'd41 )  ;
assign n3018____DOLLAR__7642 =  ( oc8051_ROM_rdata_0 ) == ( 8'd40 )  ;
assign n3019____DOLLAR__7646 =  ( oc8051_ROM_rdata_0 ) == ( 8'd39 )  ;
assign n3020____DOLLAR__7650 =  ( oc8051_ROM_rdata_0 ) == ( 8'd38 )  ;
assign n3021____DOLLAR__7654 =  ( oc8051_ROM_rdata_0 ) == ( 8'd37 )  ;
assign n3022____DOLLAR__7658 =  ( oc8051_ROM_rdata_0 ) == ( 8'd36 )  ;
assign n3023____DOLLAR__7662 =  ( oc8051_ROM_rdata_0 ) == ( 8'd35 )  ;
assign n3024____DOLLAR__7666 =  ( oc8051_ROM_rdata_0 ) == ( 8'd34 )  ;
assign n3025____DOLLAR__7670 =  ( oc8051_ROM_rdata_0 ) == ( 8'd33 )  ;
assign n3026____DOLLAR__7674 =  ( oc8051_ROM_rdata_0 ) == ( 8'd32 )  ;
assign n3027____DOLLAR__7678 =  ( oc8051_ROM_rdata_0 ) == ( 8'd31 )  ;
assign n3028____DOLLAR__7682 =  ( oc8051_ROM_rdata_0 ) == ( 8'd30 )  ;
assign n3029____DOLLAR__7686 =  ( oc8051_ROM_rdata_0 ) == ( 8'd29 )  ;
assign n3030____DOLLAR__7690 =  ( oc8051_ROM_rdata_0 ) == ( 8'd28 )  ;
assign n3031____DOLLAR__7694 =  ( oc8051_ROM_rdata_0 ) == ( 8'd27 )  ;
assign n3032____DOLLAR__7698 =  ( oc8051_ROM_rdata_0 ) == ( 8'd26 )  ;
assign n3033____DOLLAR__7702 =  ( oc8051_ROM_rdata_0 ) == ( 8'd25 )  ;
assign n3034____DOLLAR__7706 =  ( oc8051_ROM_rdata_0 ) == ( 8'd24 )  ;
assign n3035____DOLLAR__7710 =  ( oc8051_ROM_rdata_0 ) == ( 8'd23 )  ;
assign n3036____DOLLAR__7714 =  ( oc8051_ROM_rdata_0 ) == ( 8'd22 )  ;
assign n3037____DOLLAR__7718 =  ( oc8051_ROM_rdata_0 ) == ( 8'd21 )  ;
assign n3038____DOLLAR__7722 =  ( oc8051_ROM_rdata_0 ) == ( 8'd20 )  ;
assign n3039____DOLLAR__7726 =  ( oc8051_ROM_rdata_0 ) == ( 8'd19 )  ;
assign n3040____DOLLAR__7730 =  ( oc8051_ROM_rdata_0 ) == ( 8'd18 )  ;
assign n3041____DOLLAR__7734 =  ( oc8051_ROM_rdata_0 ) == ( 8'd17 )  ;
assign n3042____DOLLAR__7738 =  ( oc8051_ROM_rdata_0 ) == ( 8'd16 )  ;
assign n3043____DOLLAR__7742 =  ( oc8051_ROM_rdata_0 ) == ( 8'd15 )  ;
assign n3044____DOLLAR__7746 =  ( oc8051_ROM_rdata_0 ) == ( 8'd14 )  ;
assign n3045____DOLLAR__7750 =  ( oc8051_ROM_rdata_0 ) == ( 8'd13 )  ;
assign n3046____DOLLAR__7754 =  ( oc8051_ROM_rdata_0 ) == ( 8'd12 )  ;
assign n3047____DOLLAR__7758 =  ( oc8051_ROM_rdata_0 ) == ( 8'd11 )  ;
assign n3048____DOLLAR__7762 =  ( oc8051_ROM_rdata_0 ) == ( 8'd10 )  ;
assign n3049____DOLLAR__7766 =  ( oc8051_ROM_rdata_0 ) == ( 8'd9 )  ;
assign n3050____DOLLAR__7770 =  ( oc8051_ROM_rdata_0 ) == ( 8'd8 )  ;
assign n3051____DOLLAR__7774 =  ( oc8051_ROM_rdata_0 ) == ( 8'd7 )  ;
assign n3052____DOLLAR__7778 =  ( oc8051_ROM_rdata_0 ) == ( 8'd6 )  ;
assign n3053____DOLLAR__7782 =  ( oc8051_ROM_rdata_0 ) == ( 8'd5 )  ;
assign n3054____DOLLAR__7786 =  ( oc8051_ROM_rdata_0 ) == ( 8'd4 )  ;
assign n3055____DOLLAR__7790 =  ( oc8051_ROM_rdata_0 ) == ( 8'd3 )  ;
assign n3056____DOLLAR__7794 =  ( oc8051_ROM_rdata_0 ) == ( 8'd2 )  ;
assign n3057____DOLLAR__7798 =  ( oc8051_ROM_rdata_0 ) == ( 8'd1 )  ;
assign n3058____DOLLAR__7800 =  ( oc8051_ROM_rdata_0 ) == ( 8'd0 )  ;
assign n3059____DOLLAR__7802 =  ( n3057____DOLLAR__7798 ) | ( n3058____DOLLAR__7800 )  ;
assign n3060____DOLLAR__7803 =  ( n3056____DOLLAR__7794 ) | ( n3059____DOLLAR__7802 )  ;
assign n3061____DOLLAR__7804 =  ( n3055____DOLLAR__7790 ) | ( n3060____DOLLAR__7803 )  ;
assign n3062____DOLLAR__7805 =  ( n3054____DOLLAR__7786 ) | ( n3061____DOLLAR__7804 )  ;
assign n3063____DOLLAR__7806 =  ( n3053____DOLLAR__7782 ) | ( n3062____DOLLAR__7805 )  ;
assign n3064____DOLLAR__7807 =  ( n3052____DOLLAR__7778 ) | ( n3063____DOLLAR__7806 )  ;
assign n3065____DOLLAR__7808 =  ( n3051____DOLLAR__7774 ) | ( n3064____DOLLAR__7807 )  ;
assign n3066____DOLLAR__7809 =  ( n3050____DOLLAR__7770 ) | ( n3065____DOLLAR__7808 )  ;
assign n3067____DOLLAR__7810 =  ( n3049____DOLLAR__7766 ) | ( n3066____DOLLAR__7809 )  ;
assign n3068____DOLLAR__7811 =  ( n3048____DOLLAR__7762 ) | ( n3067____DOLLAR__7810 )  ;
assign n3069____DOLLAR__7812 =  ( n3047____DOLLAR__7758 ) | ( n3068____DOLLAR__7811 )  ;
assign n3070____DOLLAR__7813 =  ( n3046____DOLLAR__7754 ) | ( n3069____DOLLAR__7812 )  ;
assign n3071____DOLLAR__7814 =  ( n3045____DOLLAR__7750 ) | ( n3070____DOLLAR__7813 )  ;
assign n3072____DOLLAR__7815 =  ( n3044____DOLLAR__7746 ) | ( n3071____DOLLAR__7814 )  ;
assign n3073____DOLLAR__7816 =  ( n3043____DOLLAR__7742 ) | ( n3072____DOLLAR__7815 )  ;
assign n3074____DOLLAR__7817 =  ( n3042____DOLLAR__7738 ) | ( n3073____DOLLAR__7816 )  ;
assign n3075____DOLLAR__7818 =  ( n3041____DOLLAR__7734 ) | ( n3074____DOLLAR__7817 )  ;
assign n3076____DOLLAR__7819 =  ( n3040____DOLLAR__7730 ) | ( n3075____DOLLAR__7818 )  ;
assign n3077____DOLLAR__7820 =  ( n3039____DOLLAR__7726 ) | ( n3076____DOLLAR__7819 )  ;
assign n3078____DOLLAR__7821 =  ( n3038____DOLLAR__7722 ) | ( n3077____DOLLAR__7820 )  ;
assign n3079____DOLLAR__7822 =  ( n3037____DOLLAR__7718 ) | ( n3078____DOLLAR__7821 )  ;
assign n3080____DOLLAR__7823 =  ( n3036____DOLLAR__7714 ) | ( n3079____DOLLAR__7822 )  ;
assign n3081____DOLLAR__7824 =  ( n3035____DOLLAR__7710 ) | ( n3080____DOLLAR__7823 )  ;
assign n3082____DOLLAR__7825 =  ( n3034____DOLLAR__7706 ) | ( n3081____DOLLAR__7824 )  ;
assign n3083____DOLLAR__7826 =  ( n3033____DOLLAR__7702 ) | ( n3082____DOLLAR__7825 )  ;
assign n3084____DOLLAR__7827 =  ( n3032____DOLLAR__7698 ) | ( n3083____DOLLAR__7826 )  ;
assign n3085____DOLLAR__7828 =  ( n3031____DOLLAR__7694 ) | ( n3084____DOLLAR__7827 )  ;
assign n3086____DOLLAR__7829 =  ( n3030____DOLLAR__7690 ) | ( n3085____DOLLAR__7828 )  ;
assign n3087____DOLLAR__7830 =  ( n3029____DOLLAR__7686 ) | ( n3086____DOLLAR__7829 )  ;
assign n3088____DOLLAR__7831 =  ( n3028____DOLLAR__7682 ) | ( n3087____DOLLAR__7830 )  ;
assign n3089____DOLLAR__7832 =  ( n3027____DOLLAR__7678 ) | ( n3088____DOLLAR__7831 )  ;
assign n3090____DOLLAR__7833 =  ( n3026____DOLLAR__7674 ) | ( n3089____DOLLAR__7832 )  ;
assign n3091____DOLLAR__7834 =  ( n3025____DOLLAR__7670 ) | ( n3090____DOLLAR__7833 )  ;
assign n3092____DOLLAR__7835 =  ( n3024____DOLLAR__7666 ) | ( n3091____DOLLAR__7834 )  ;
assign n3093____DOLLAR__7836 =  ( n3023____DOLLAR__7662 ) | ( n3092____DOLLAR__7835 )  ;
assign n3094____DOLLAR__7837 =  ( n3022____DOLLAR__7658 ) | ( n3093____DOLLAR__7836 )  ;
assign n3095____DOLLAR__7838 =  ( n3021____DOLLAR__7654 ) | ( n3094____DOLLAR__7837 )  ;
assign n3096____DOLLAR__7839 =  ( n3020____DOLLAR__7650 ) | ( n3095____DOLLAR__7838 )  ;
assign n3097____DOLLAR__7840 =  ( n3019____DOLLAR__7646 ) | ( n3096____DOLLAR__7839 )  ;
assign n3098____DOLLAR__7841 =  ( n3018____DOLLAR__7642 ) | ( n3097____DOLLAR__7840 )  ;
assign n3099____DOLLAR__7842 =  ( n3017____DOLLAR__7638 ) | ( n3098____DOLLAR__7841 )  ;
assign n3100____DOLLAR__7843 =  ( n3016____DOLLAR__7634 ) | ( n3099____DOLLAR__7842 )  ;
assign n3101____DOLLAR__7844 =  ( n3015____DOLLAR__7630 ) | ( n3100____DOLLAR__7843 )  ;
assign n3102____DOLLAR__7845 =  ( n3014____DOLLAR__7626 ) | ( n3101____DOLLAR__7844 )  ;
assign n3103____DOLLAR__7846 =  ( n3013____DOLLAR__7622 ) | ( n3102____DOLLAR__7845 )  ;
assign n3104____DOLLAR__7847 =  ( n3012____DOLLAR__7618 ) | ( n3103____DOLLAR__7846 )  ;
assign n3105____DOLLAR__7848 =  ( n3011____DOLLAR__7614 ) | ( n3104____DOLLAR__7847 )  ;
assign n3106____DOLLAR__7849 =  ( n3010____DOLLAR__7610 ) | ( n3105____DOLLAR__7848 )  ;
assign n3107____DOLLAR__7850 =  ( n3009____DOLLAR__7606 ) | ( n3106____DOLLAR__7849 )  ;
assign n3108____DOLLAR__7851 =  ( n3008____DOLLAR__7602 ) | ( n3107____DOLLAR__7850 )  ;
assign n3109____DOLLAR__7852 =  ( n3007____DOLLAR__7598 ) | ( n3108____DOLLAR__7851 )  ;
assign n3110____DOLLAR__7853 =  ( n3006____DOLLAR__7594 ) | ( n3109____DOLLAR__7852 )  ;
assign n3111____DOLLAR__7854 =  ( n3005____DOLLAR__7590 ) | ( n3110____DOLLAR__7853 )  ;
assign n3112____DOLLAR__7855 =  ( n3004____DOLLAR__7586 ) | ( n3111____DOLLAR__7854 )  ;
assign n3113____DOLLAR__7856 =  ( n3003____DOLLAR__7582 ) | ( n3112____DOLLAR__7855 )  ;
assign n3114____DOLLAR__7857 =  ( n3002____DOLLAR__7578 ) | ( n3113____DOLLAR__7856 )  ;
assign n3115____DOLLAR__7858 =  ( n3001____DOLLAR__7574 ) | ( n3114____DOLLAR__7857 )  ;
assign n3116____DOLLAR__7859 =  ( n3000____DOLLAR__7570 ) | ( n3115____DOLLAR__7858 )  ;
assign n3117____DOLLAR__7860 =  ( n2999____DOLLAR__7566 ) | ( n3116____DOLLAR__7859 )  ;
assign n3118____DOLLAR__7861 =  ( n2998____DOLLAR__7562 ) | ( n3117____DOLLAR__7860 )  ;
assign n3119____DOLLAR__7862 =  ( n2997____DOLLAR__7558 ) | ( n3118____DOLLAR__7861 )  ;
assign n3120____DOLLAR__7863 =  ( n2996____DOLLAR__7554 ) | ( n3119____DOLLAR__7862 )  ;
assign n3121____DOLLAR__7864 =  ( n2995____DOLLAR__7550 ) | ( n3120____DOLLAR__7863 )  ;
assign n3122____DOLLAR__7865 =  ( n2994____DOLLAR__7546 ) | ( n3121____DOLLAR__7864 )  ;
assign n3123____DOLLAR__7866 =  ( n2993____DOLLAR__7542 ) | ( n3122____DOLLAR__7865 )  ;
assign n3124____DOLLAR__7867 =  ( n2992____DOLLAR__7538 ) | ( n3123____DOLLAR__7866 )  ;
assign n3125____DOLLAR__7868 =  ( n2991____DOLLAR__7534 ) | ( n3124____DOLLAR__7867 )  ;
assign n3126____DOLLAR__7869 =  ( n2990____DOLLAR__7530 ) | ( n3125____DOLLAR__7868 )  ;
assign n3127____DOLLAR__7870 =  ( n2989____DOLLAR__7526 ) | ( n3126____DOLLAR__7869 )  ;
assign n3128____DOLLAR__7871 =  ( n2988____DOLLAR__7522 ) | ( n3127____DOLLAR__7870 )  ;
assign n3129____DOLLAR__7872 =  ( n2987____DOLLAR__7518 ) | ( n3128____DOLLAR__7871 )  ;
assign n3130____DOLLAR__7873 =  ( n2986____DOLLAR__7514 ) | ( n3129____DOLLAR__7872 )  ;
assign n3131____DOLLAR__7874 =  ( n2985____DOLLAR__7510 ) | ( n3130____DOLLAR__7873 )  ;
assign n3132____DOLLAR__7875 =  ( n2984____DOLLAR__7506 ) | ( n3131____DOLLAR__7874 )  ;
assign n3133____DOLLAR__7876 =  ( n2983____DOLLAR__7502 ) | ( n3132____DOLLAR__7875 )  ;
assign n3134____DOLLAR__7877 =  ( n2982____DOLLAR__7498 ) | ( n3133____DOLLAR__7876 )  ;
assign n3135____DOLLAR__7878 =  ( n2981____DOLLAR__7494 ) | ( n3134____DOLLAR__7877 )  ;
assign n3136____DOLLAR__7879 =  ( n2980____DOLLAR__7490 ) | ( n3135____DOLLAR__7878 )  ;
assign n3137____DOLLAR__7880 =  ( n2979____DOLLAR__7486 ) | ( n3136____DOLLAR__7879 )  ;
assign n3138____DOLLAR__7881 =  ( n2978____DOLLAR__7482 ) | ( n3137____DOLLAR__7880 )  ;
assign n3139____DOLLAR__7882 =  ( n2977____DOLLAR__7478 ) | ( n3138____DOLLAR__7881 )  ;
assign n3140____DOLLAR__7883 =  ( n2976____DOLLAR__7474 ) | ( n3139____DOLLAR__7882 )  ;
assign n3141____DOLLAR__7884 =  ( n2975____DOLLAR__7470 ) | ( n3140____DOLLAR__7883 )  ;
assign n3142____DOLLAR__7885 =  ( n2974____DOLLAR__7466 ) | ( n3141____DOLLAR__7884 )  ;
assign n3143____DOLLAR__7886 =  ( n2973____DOLLAR__7462 ) | ( n3142____DOLLAR__7885 )  ;
assign n3144____DOLLAR__7887 =  ( n2972____DOLLAR__7458 ) | ( n3143____DOLLAR__7886 )  ;
assign n3145____DOLLAR__7888 =  ( n2971____DOLLAR__7454 ) | ( n3144____DOLLAR__7887 )  ;
assign n3146____DOLLAR__7889 =  ( n2970____DOLLAR__7450 ) | ( n3145____DOLLAR__7888 )  ;
assign n3147____DOLLAR__7890 =  ( n2969____DOLLAR__7446 ) | ( n3146____DOLLAR__7889 )  ;
assign n3148____DOLLAR__7891 =  ( n2968____DOLLAR__7442 ) | ( n3147____DOLLAR__7890 )  ;
assign n3149____DOLLAR__7892 =  ( n2967____DOLLAR__7438 ) | ( n3148____DOLLAR__7891 )  ;
assign n3150____DOLLAR__7893 =  ( n2966____DOLLAR__7434 ) | ( n3149____DOLLAR__7892 )  ;
assign n3151____DOLLAR__7894 =  ( n2965____DOLLAR__7430 ) | ( n3150____DOLLAR__7893 )  ;
assign n3152____DOLLAR__7895 =  ( n2964____DOLLAR__7426 ) | ( n3151____DOLLAR__7894 )  ;
assign n3153____DOLLAR__7896 =  ( n2963____DOLLAR__7422 ) | ( n3152____DOLLAR__7895 )  ;
assign n3154____DOLLAR__7897 =  ( n2962____DOLLAR__7418 ) | ( n3153____DOLLAR__7896 )  ;
assign n3155____DOLLAR__7898 =  ( n2961____DOLLAR__7414 ) | ( n3154____DOLLAR__7897 )  ;
assign n3156____DOLLAR__7899 =  ( n2960____DOLLAR__7410 ) | ( n3155____DOLLAR__7898 )  ;
assign n3157____DOLLAR__7900 =  ( n2959____DOLLAR__7406 ) | ( n3156____DOLLAR__7899 )  ;
assign n3158____DOLLAR__7901 =  ( n2958____DOLLAR__7402 ) | ( n3157____DOLLAR__7900 )  ;
assign n3159____DOLLAR__7902 =  ( n2957____DOLLAR__7398 ) | ( n3158____DOLLAR__7901 )  ;
assign n3160____DOLLAR__7903 =  ( n2956____DOLLAR__7394 ) | ( n3159____DOLLAR__7902 )  ;
assign n3161____DOLLAR__7904 =  ( n2955____DOLLAR__7390 ) | ( n3160____DOLLAR__7903 )  ;
assign n3162____DOLLAR__7905 =  ( n2954____DOLLAR__7386 ) | ( n3161____DOLLAR__7904 )  ;
assign n3163____DOLLAR__7906 =  ( n2953____DOLLAR__7382 ) | ( n3162____DOLLAR__7905 )  ;
assign n3164____DOLLAR__7907 =  ( n2952____DOLLAR__7378 ) | ( n3163____DOLLAR__7906 )  ;
assign n3165____DOLLAR__7908 =  ( n2951____DOLLAR__7374 ) | ( n3164____DOLLAR__7907 )  ;
assign n3166____DOLLAR__7909 =  ( n2950____DOLLAR__7370 ) | ( n3165____DOLLAR__7908 )  ;
assign n3167____DOLLAR__7910 =  ( n2949____DOLLAR__7366 ) | ( n3166____DOLLAR__7909 )  ;
assign n3168____DOLLAR__7911 =  ( n2948____DOLLAR__7362 ) | ( n3167____DOLLAR__7910 )  ;
assign n3169____DOLLAR__7912 =  ( n2947____DOLLAR__7358 ) | ( n3168____DOLLAR__7911 )  ;
assign n3170____DOLLAR__7913 =  ( n2946____DOLLAR__7354 ) | ( n3169____DOLLAR__7912 )  ;
assign n3171____DOLLAR__7914 =  ( n2945____DOLLAR__7350 ) | ( n3170____DOLLAR__7913 )  ;
assign n3172____DOLLAR__7915 =  ( n2944____DOLLAR__7346 ) | ( n3171____DOLLAR__7914 )  ;
assign n3173____DOLLAR__7916 =  ( n2943____DOLLAR__7342 ) | ( n3172____DOLLAR__7915 )  ;
assign n3174____DOLLAR__7917 =  ( n2942____DOLLAR__7338 ) | ( n3173____DOLLAR__7916 )  ;
assign n3175____DOLLAR__7918 =  ( n2941____DOLLAR__7334 ) | ( n3174____DOLLAR__7917 )  ;
assign n3176____DOLLAR__7919 =  ( n2940____DOLLAR__7330 ) | ( n3175____DOLLAR__7918 )  ;
assign n3177____DOLLAR__7920 =  ( n2939____DOLLAR__7326 ) | ( n3176____DOLLAR__7919 )  ;
assign n3178____DOLLAR__7921 =  ( n2938____DOLLAR__7322 ) | ( n3177____DOLLAR__7920 )  ;
assign n3179____DOLLAR__7922 =  ( n2937____DOLLAR__7318 ) | ( n3178____DOLLAR__7921 )  ;
assign n3180____DOLLAR__7923 =  ( n2936____DOLLAR__7314 ) | ( n3179____DOLLAR__7922 )  ;
assign n3181____DOLLAR__7924 =  ( n2935____DOLLAR__7310 ) | ( n3180____DOLLAR__7923 )  ;
assign n3182____DOLLAR__7925 =  ( n2934____DOLLAR__7306 ) | ( n3181____DOLLAR__7924 )  ;
assign n3183____DOLLAR__7926 =  ( n2933____DOLLAR__7302 ) | ( n3182____DOLLAR__7925 )  ;
assign n3184____DOLLAR__7927 =  ( n2932____DOLLAR__7298 ) | ( n3183____DOLLAR__7926 )  ;
assign n3185____DOLLAR__7928 =  ( n2931____DOLLAR__7294 ) | ( n3184____DOLLAR__7927 )  ;
assign n3186____DOLLAR__7929 =  ( n2930____DOLLAR__7290 ) | ( n3185____DOLLAR__7928 )  ;
assign n3187____DOLLAR__7930 =  ( n2929____DOLLAR__7286 ) | ( n3186____DOLLAR__7929 )  ;
assign n3188____DOLLAR__7931 =  ( n2928____DOLLAR__7282 ) | ( n3187____DOLLAR__7930 )  ;
assign n3189____DOLLAR__7932 =  ( n2927____DOLLAR__7278 ) | ( n3188____DOLLAR__7931 )  ;
assign n3190____DOLLAR__7933 =  ( n2926____DOLLAR__7274 ) | ( n3189____DOLLAR__7932 )  ;
assign n3191____DOLLAR__7934 =  ( n2925____DOLLAR__7270 ) | ( n3190____DOLLAR__7933 )  ;
assign n3192____DOLLAR__7935 =  ( n2924____DOLLAR__7266 ) | ( n3191____DOLLAR__7934 )  ;
assign n3193____DOLLAR__7936 =  ( n2923____DOLLAR__7262 ) | ( n3192____DOLLAR__7935 )  ;
assign n3194____DOLLAR__7937 =  ( n2922____DOLLAR__7258 ) | ( n3193____DOLLAR__7936 )  ;
assign n3195____DOLLAR__7938 =  ( n2921____DOLLAR__7254 ) | ( n3194____DOLLAR__7937 )  ;
assign n3196____DOLLAR__7939 =  ( n2920____DOLLAR__7250 ) | ( n3195____DOLLAR__7938 )  ;
assign n3197____DOLLAR__7940 =  ( n2919____DOLLAR__7246 ) | ( n3196____DOLLAR__7939 )  ;
assign n3198____DOLLAR__7941 =  ( n2918____DOLLAR__7242 ) | ( n3197____DOLLAR__7940 )  ;
assign n3199____DOLLAR__7942 =  ( n2917____DOLLAR__7238 ) | ( n3198____DOLLAR__7941 )  ;
assign n3200____DOLLAR__7943 =  ( n2916____DOLLAR__7234 ) | ( n3199____DOLLAR__7942 )  ;
assign n3201____DOLLAR__7944 =  ( n2915____DOLLAR__7230 ) | ( n3200____DOLLAR__7943 )  ;
assign n3202____DOLLAR__7945 =  ( n2914____DOLLAR__7226 ) | ( n3201____DOLLAR__7944 )  ;
assign n3203____DOLLAR__7946 =  ( n2913____DOLLAR__7222 ) | ( n3202____DOLLAR__7945 )  ;
assign n3204____DOLLAR__7947 =  ( n2912____DOLLAR__7218 ) | ( n3203____DOLLAR__7946 )  ;
assign n3205____DOLLAR__7948 =  ( n2911____DOLLAR__7214 ) | ( n3204____DOLLAR__7947 )  ;
assign n3206____DOLLAR__7949 =  ( n2910____DOLLAR__7210 ) | ( n3205____DOLLAR__7948 )  ;
assign n3207____DOLLAR__7950 =  ( n2909____DOLLAR__7206 ) | ( n3206____DOLLAR__7949 )  ;
assign n3208____DOLLAR__7951 =  ( n2908____DOLLAR__7202 ) | ( n3207____DOLLAR__7950 )  ;
assign n3209____DOLLAR__7952 =  ( n2907____DOLLAR__7198 ) | ( n3208____DOLLAR__7951 )  ;
assign n3210____DOLLAR__7953 =  ( n2906____DOLLAR__7194 ) | ( n3209____DOLLAR__7952 )  ;
assign n3211____DOLLAR__7954 =  ( n2905____DOLLAR__7190 ) | ( n3210____DOLLAR__7953 )  ;
assign n3212____DOLLAR__7955 =  ( n2904____DOLLAR__7186 ) | ( n3211____DOLLAR__7954 )  ;
assign n3213____DOLLAR__7956 =  ( n2903____DOLLAR__7182 ) | ( n3212____DOLLAR__7955 )  ;
assign n3214____DOLLAR__7957 =  ( n2902____DOLLAR__7178 ) | ( n3213____DOLLAR__7956 )  ;
assign n3215____DOLLAR__7958 =  ( n2901____DOLLAR__7174 ) | ( n3214____DOLLAR__7957 )  ;
assign n3216____DOLLAR__7959 =  ( n2900____DOLLAR__7170 ) | ( n3215____DOLLAR__7958 )  ;
assign n3217____DOLLAR__7960 =  ( n2899____DOLLAR__7166 ) | ( n3216____DOLLAR__7959 )  ;
assign n3218____DOLLAR__7961 =  ( n2898____DOLLAR__7162 ) | ( n3217____DOLLAR__7960 )  ;
assign n3219____DOLLAR__7962 =  ( n2897____DOLLAR__7158 ) | ( n3218____DOLLAR__7961 )  ;
assign n3220____DOLLAR__7963 =  ( n2896____DOLLAR__7154 ) | ( n3219____DOLLAR__7962 )  ;
assign n3221____DOLLAR__7964 =  ( n2895____DOLLAR__7150 ) | ( n3220____DOLLAR__7963 )  ;
assign n3222____DOLLAR__7965 =  ( n2894____DOLLAR__7146 ) | ( n3221____DOLLAR__7964 )  ;
assign n3223____DOLLAR__7966 =  ( n2893____DOLLAR__7142 ) | ( n3222____DOLLAR__7965 )  ;
assign n3224____DOLLAR__7967 =  ( n2892____DOLLAR__7138 ) | ( n3223____DOLLAR__7966 )  ;
assign n3225____DOLLAR__7968 =  ( n2891____DOLLAR__7134 ) | ( n3224____DOLLAR__7967 )  ;
assign n3226____DOLLAR__7969 =  ( n2890____DOLLAR__7130 ) | ( n3225____DOLLAR__7968 )  ;
assign n3227____DOLLAR__7970 =  ( n2889____DOLLAR__7126 ) | ( n3226____DOLLAR__7969 )  ;
assign n3228____DOLLAR__7971 =  ( n2888____DOLLAR__7122 ) | ( n3227____DOLLAR__7970 )  ;
assign n3229____DOLLAR__7972 =  ( n2887____DOLLAR__7118 ) | ( n3228____DOLLAR__7971 )  ;
assign n3230____DOLLAR__7973 =  ( n2886____DOLLAR__7114 ) | ( n3229____DOLLAR__7972 )  ;
assign n3231____DOLLAR__7974 =  ( n2885____DOLLAR__7110 ) | ( n3230____DOLLAR__7973 )  ;
assign n3232____DOLLAR__7975 =  ( n2884____DOLLAR__7106 ) | ( n3231____DOLLAR__7974 )  ;
assign n3233____DOLLAR__7976 =  ( n2883____DOLLAR__7102 ) | ( n3232____DOLLAR__7975 )  ;
assign n3234____DOLLAR__7977 =  ( n2882____DOLLAR__7098 ) | ( n3233____DOLLAR__7976 )  ;
assign n3235____DOLLAR__7978 =  ( n2881____DOLLAR__7094 ) | ( n3234____DOLLAR__7977 )  ;
assign n3236____DOLLAR__7979 =  ( n2880____DOLLAR__7090 ) | ( n3235____DOLLAR__7978 )  ;
assign n3237____DOLLAR__7980 =  ( n2879____DOLLAR__7086 ) | ( n3236____DOLLAR__7979 )  ;
assign n3238____DOLLAR__7981 =  ( n2878____DOLLAR__7082 ) | ( n3237____DOLLAR__7980 )  ;
assign n3239____DOLLAR__7982 =  ( n2877____DOLLAR__7078 ) | ( n3238____DOLLAR__7981 )  ;
assign n3240____DOLLAR__7983 =  ( n2876____DOLLAR__7074 ) | ( n3239____DOLLAR__7982 )  ;
assign n3241____DOLLAR__7984 =  ( n2875____DOLLAR__7070 ) | ( n3240____DOLLAR__7983 )  ;
assign n3242____DOLLAR__7985 =  ( n2874____DOLLAR__7066 ) | ( n3241____DOLLAR__7984 )  ;
assign n3243____DOLLAR__7986 =  ( n2873____DOLLAR__7062 ) | ( n3242____DOLLAR__7985 )  ;
assign n3244____DOLLAR__7987 =  ( n2872____DOLLAR__7058 ) | ( n3243____DOLLAR__7986 )  ;
assign n3245____DOLLAR__7988 =  ( n2871____DOLLAR__7054 ) | ( n3244____DOLLAR__7987 )  ;
assign n3246____DOLLAR__7989 =  ( n2870____DOLLAR__7050 ) | ( n3245____DOLLAR__7988 )  ;
assign n3247____DOLLAR__7990 =  ( n2869____DOLLAR__7046 ) | ( n3246____DOLLAR__7989 )  ;
assign n3248____DOLLAR__7991 =  ( n2868____DOLLAR__7042 ) | ( n3247____DOLLAR__7990 )  ;
assign n3249____DOLLAR__7992 =  ( n2867____DOLLAR__7038 ) | ( n3248____DOLLAR__7991 )  ;
assign n3250____DOLLAR__7993 =  ( n2866____DOLLAR__7034 ) | ( n3249____DOLLAR__7992 )  ;
assign n3251____DOLLAR__7994 =  ( n2865____DOLLAR__7030 ) | ( n3250____DOLLAR__7993 )  ;
assign n3252____DOLLAR__7995 =  ( n2864____DOLLAR__7026 ) | ( n3251____DOLLAR__7994 )  ;
assign n3253____DOLLAR__7996 =  ( n2863____DOLLAR__7022 ) | ( n3252____DOLLAR__7995 )  ;
assign n3254____DOLLAR__7997 =  ( n2862____DOLLAR__7018 ) | ( n3253____DOLLAR__7996 )  ;
assign n3255____DOLLAR__7998 =  ( n2861____DOLLAR__7014 ) | ( n3254____DOLLAR__7997 )  ;
assign n3256____DOLLAR__7999 =  ( n2860____DOLLAR__7010 ) | ( n3255____DOLLAR__7998 )  ;
assign n3257____DOLLAR__8000 =  ( n2859____DOLLAR__7006 ) | ( n3256____DOLLAR__7999 )  ;
assign n3258____DOLLAR__8001 =  ( n2858____DOLLAR__7002 ) | ( n3257____DOLLAR__8000 )  ;
assign n3259____DOLLAR__8002 =  ( n2857____DOLLAR__6998 ) | ( n3258____DOLLAR__8001 )  ;
assign n3260____DOLLAR__8003 =  ( n2856____DOLLAR__6994 ) | ( n3259____DOLLAR__8002 )  ;
assign n3261____DOLLAR__8004 =  ( n2855____DOLLAR__6990 ) | ( n3260____DOLLAR__8003 )  ;
assign n3262____DOLLAR__8005 =  ( n2854____DOLLAR__6986 ) | ( n3261____DOLLAR__8004 )  ;
assign n3263____DOLLAR__8006 =  ( n2853____DOLLAR__6982 ) | ( n3262____DOLLAR__8005 )  ;
assign n3264____DOLLAR__8007 =  ( n2852____DOLLAR__6978 ) | ( n3263____DOLLAR__8006 )  ;
assign n3265____DOLLAR__8008 =  ( n2851____DOLLAR__6974 ) | ( n3264____DOLLAR__8007 )  ;
assign n3266____DOLLAR__8009 =  ( n2850____DOLLAR__6970 ) | ( n3265____DOLLAR__8008 )  ;
assign n3267____DOLLAR__8010 =  ( n2849____DOLLAR__6966 ) | ( n3266____DOLLAR__8009 )  ;
assign n3268____DOLLAR__8011 =  ( n2848____DOLLAR__6962 ) | ( n3267____DOLLAR__8010 )  ;
assign n3269____DOLLAR__8012 =  ( n2847____DOLLAR__6958 ) | ( n3268____DOLLAR__8011 )  ;
assign n3270____DOLLAR__8013 =  ( n2846____DOLLAR__6954 ) | ( n3269____DOLLAR__8012 )  ;
assign n3271____DOLLAR__8014 =  ( n2845____DOLLAR__6950 ) | ( n3270____DOLLAR__8013 )  ;
assign n3272____DOLLAR__8015 =  ( n2844____DOLLAR__6946 ) | ( n3271____DOLLAR__8014 )  ;
assign n3273____DOLLAR__8016 =  ( n2843____DOLLAR__6942 ) | ( n3272____DOLLAR__8015 )  ;
assign n3274____DOLLAR__8017 =  ( n2842____DOLLAR__6938 ) | ( n3273____DOLLAR__8016 )  ;
assign n3275____DOLLAR__8018 =  ( n2841____DOLLAR__6934 ) | ( n3274____DOLLAR__8017 )  ;
assign n3276____DOLLAR__8019 =  ( n2840____DOLLAR__6930 ) | ( n3275____DOLLAR__8018 )  ;
assign n3277____DOLLAR__8020 =  ( n2839____DOLLAR__6926 ) | ( n3276____DOLLAR__8019 )  ;
assign n3278____DOLLAR__8021 =  ( n2838____DOLLAR__6922 ) | ( n3277____DOLLAR__8020 )  ;
assign n3279____DOLLAR__8022 =  ( n2837____DOLLAR__6918 ) | ( n3278____DOLLAR__8021 )  ;
assign n3280____DOLLAR__8023 =  ( n2836____DOLLAR__6914 ) | ( n3279____DOLLAR__8022 )  ;
assign n3281____DOLLAR__8024 =  ( n2835____DOLLAR__6910 ) | ( n3280____DOLLAR__8023 )  ;
assign n3282____DOLLAR__8025 =  ( n2834____DOLLAR__6906 ) | ( n3281____DOLLAR__8024 )  ;
assign n3283____DOLLAR__8026 =  ( n2833____DOLLAR__6902 ) | ( n3282____DOLLAR__8025 )  ;
assign n3284____DOLLAR__8027 =  ( n2832____DOLLAR__6898 ) | ( n3283____DOLLAR__8026 )  ;
assign n3285____DOLLAR__8028 =  ( n2831____DOLLAR__6894 ) | ( n3284____DOLLAR__8027 )  ;
assign n3286____DOLLAR__8029 =  ( n2830____DOLLAR__6890 ) | ( n3285____DOLLAR__8028 )  ;
assign n3287____DOLLAR__8030 =  ( n2829____DOLLAR__6886 ) | ( n3286____DOLLAR__8029 )  ;
assign n3288____DOLLAR__8031 =  ( n2828____DOLLAR__6882 ) | ( n3287____DOLLAR__8030 )  ;
assign n3289____DOLLAR__8032 =  ( n2827____DOLLAR__6878 ) | ( n3288____DOLLAR__8031 )  ;
assign n3290____DOLLAR__8033 =  ( n2826____DOLLAR__6874 ) | ( n3289____DOLLAR__8032 )  ;
assign n3291____DOLLAR__8034 =  ( n2825____DOLLAR__6870 ) | ( n3290____DOLLAR__8033 )  ;
assign n3292____DOLLAR__8035 =  ( n2824____DOLLAR__6866 ) | ( n3291____DOLLAR__8034 )  ;
assign n3293____DOLLAR__8036 =  ( n2823____DOLLAR__6862 ) | ( n3292____DOLLAR__8035 )  ;
assign n3294____DOLLAR__8037 =  ( n2822____DOLLAR__6858 ) | ( n3293____DOLLAR__8036 )  ;
assign n3295____DOLLAR__8038 =  ( n2821____DOLLAR__6854 ) | ( n3294____DOLLAR__8037 )  ;
assign n3296____DOLLAR__8039 =  ( n2820____DOLLAR__6850 ) | ( n3295____DOLLAR__8038 )  ;
assign n3297____DOLLAR__8040 =  ( n2819____DOLLAR__6846 ) | ( n3296____DOLLAR__8039 )  ;
assign n3298____DOLLAR__8041 =  ( n2818____DOLLAR__6842 ) | ( n3297____DOLLAR__8040 )  ;
assign n3299____DOLLAR__8042 =  ( n2817____DOLLAR__6838 ) | ( n3298____DOLLAR__8041 )  ;
assign n3300____DOLLAR__8043 =  ( n2816____DOLLAR__6834 ) | ( n3299____DOLLAR__8042 )  ;
assign n3301____DOLLAR__8044 =  ( n2815____DOLLAR__6830 ) | ( n3300____DOLLAR__8043 )  ;
assign n3302____DOLLAR__8045 =  ( n2814____DOLLAR__6826 ) | ( n3301____DOLLAR__8044 )  ;
assign n3303____DOLLAR__8046 =  ( n2813____DOLLAR__6822 ) | ( n3302____DOLLAR__8045 )  ;
assign n3304____DOLLAR__8047 =  ( n2812____DOLLAR__6818 ) | ( n3303____DOLLAR__8046 )  ;
assign n3305____DOLLAR__8048 =  ( n2811____DOLLAR__6814 ) | ( n3304____DOLLAR__8047 )  ;
assign n3306____DOLLAR__8049 =  ( n2810____DOLLAR__6810 ) | ( n3305____DOLLAR__8048 )  ;
assign n3307____DOLLAR__8050 =  ( n2809____DOLLAR__6806 ) | ( n3306____DOLLAR__8049 )  ;
assign n3308____DOLLAR__8051 =  ( n2808____DOLLAR__6802 ) | ( n3307____DOLLAR__8050 )  ;
assign n3309____DOLLAR__8052 =  ( n2807____DOLLAR__6798 ) | ( n3308____DOLLAR__8051 )  ;
assign n3310____DOLLAR__8053 =  ( n2806____DOLLAR__6794 ) | ( n3309____DOLLAR__8052 )  ;
assign n3311____DOLLAR__8056 =  ( n3310____DOLLAR__8053 ) ? ( 8'd0 ) : ( XRAM_DATA_OUT ) ;
assign n3312____DOLLAR__8057 =  ( n2805____DOLLAR__6789 ) ? ( ACC ) : ( n3311____DOLLAR__8056 ) ;
assign n3313____DOLLAR__203215 =  ( PC ) + ( 16'd1 )  ;
assign n3314____DOLLAR__203218 =  ( PC ) + ( 16'd2 )  ;
assign n3315____DOLLAR__203842 =  ( aes_status ) == ( 2'd0 )  ;
assign n3316____DOLLAR__204105 = ~ ( n3315____DOLLAR__203842 )  ;
assign n3317____DOLLAR__204106 =  ( n0____DOLLAR__167758 ) & (n3316____DOLLAR__204105 )  ;
assign n3318____DOLLAR__204104 =  ( n0____DOLLAR__167758 ) & (n3315____DOLLAR__203842 )  ;
assign n3319____DOLLAR__203240 =  { ( DPH ) , ( DPL ) }  ;
assign n3320____DOLLAR__203836 =  ( n3319____DOLLAR__203240 ) < ( 16'd65280 )  ;
assign n3321____DOLLAR__203829 =  ( n3319____DOLLAR__203240 ) == ( 16'd65344 )  ;
assign n3322____DOLLAR__203831 =  ( n3319____DOLLAR__203240 ) > ( 16'd65344 )  ;
assign n3323____DOLLAR__203833 =  ( n3321____DOLLAR__203829 ) | ( n3322____DOLLAR__203831 )  ;
assign n3324____DOLLAR__203838 =  ( n3320____DOLLAR__203836 ) | ( n3323____DOLLAR__203833 )  ;
assign n3325____DOLLAR__204108 = ~ ( n3324____DOLLAR__203838 )  ;
assign n3326____DOLLAR__204109 =  ( n3318____DOLLAR__204104 ) & (n3325____DOLLAR__204108 )  ;
assign n3327____DOLLAR__204107 =  ( n3318____DOLLAR__204104 ) & (n3324____DOLLAR__203838 )  ;
assign XRAM_addr0 = n3327____DOLLAR__204107 ? (n3319____DOLLAR__203240) : (0) ;
assign XRAM_data0 = n3327____DOLLAR__204107 ? (ACC) : ('d0) ;
assign XRAM_wen0 = (n3327____DOLLAR__204107)&&__START__ ? ( 1'b1 ) : (1'b0) ;
assign n3328____DOLLAR__203301 =  ( aes_status ) == ( 2'd0 )  ;
assign n3329____DOLLAR__203296 =  ( n3319____DOLLAR__203240 ) == ( 16'd65282 )  ;
assign n3330____DOLLAR__203286 = aes_address[15:8] ;
assign n3331____DOLLAR__203292 =  { ( n3330____DOLLAR__203286 ) , ( ACC ) }  ;
assign n3332____DOLLAR__203283 =  ( n3319____DOLLAR__203240 ) == ( 16'd65283 )  ;
assign n3333____DOLLAR__203273 = aes_address[7:0] ;
assign n3334____DOLLAR__203279 =  { ( ACC ) , ( n3333____DOLLAR__203273 ) }  ;
assign n3335____DOLLAR__203285 =  ( n3332____DOLLAR__203283 ) ? ( n3334____DOLLAR__203279 ) : ( aes_address ) ;
assign n3336____DOLLAR__203298 =  ( n3329____DOLLAR__203296 ) ? ( n3331____DOLLAR__203292 ) : ( n3335____DOLLAR__203285 ) ;
assign n3337____DOLLAR__203303 =  ( n3328____DOLLAR__203301 ) ? ( n3336____DOLLAR__203298 ) : ( aes_address ) ;
assign n3338____DOLLAR__203270 =  ( aes_status ) == ( 2'd0 )  ;
assign n3339____DOLLAR__203265 =  ( n3319____DOLLAR__203240 ) == ( 16'd65284 )  ;
assign n3340____DOLLAR__203255 = aes_length[15:8] ;
assign n3341____DOLLAR__203261 =  { ( n3340____DOLLAR__203255 ) , ( ACC ) }  ;
assign n3342____DOLLAR__203252 =  ( n3319____DOLLAR__203240 ) == ( 16'd65285 )  ;
assign n3343____DOLLAR__203242 = aes_length[7:0] ;
assign n3344____DOLLAR__203248 =  { ( ACC ) , ( n3343____DOLLAR__203242 ) }  ;
assign n3345____DOLLAR__203254 =  ( n3342____DOLLAR__203252 ) ? ( n3344____DOLLAR__203248 ) : ( aes_length ) ;
assign n3346____DOLLAR__203267 =  ( n3339____DOLLAR__203265 ) ? ( n3341____DOLLAR__203261 ) : ( n3345____DOLLAR__203254 ) ;
assign n3347____DOLLAR__203272 =  ( n3338____DOLLAR__203270 ) ? ( n3346____DOLLAR__203267 ) : ( aes_length ) ;
assign n3348____DOLLAR__203556 =  ( aes_status ) == ( 2'd0 )  ;
assign n3349____DOLLAR__203542 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3350____DOLLAR__203545 =  ( n3349____DOLLAR__203542 ) == ( 16'd15 )  ;
assign n3351____DOLLAR__203538 = aes_key[127:120] ;
assign n3352____DOLLAR__203547 =  ( n3350____DOLLAR__203545 ) ? ( ACC ) : ( n3351____DOLLAR__203538 ) ;
assign n3353____DOLLAR__203526 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3354____DOLLAR__203529 =  ( n3353____DOLLAR__203526 ) == ( 16'd14 )  ;
assign n3355____DOLLAR__203522 = aes_key[119:112] ;
assign n3356____DOLLAR__203531 =  ( n3354____DOLLAR__203529 ) ? ( ACC ) : ( n3355____DOLLAR__203522 ) ;
assign n3357____DOLLAR__203510 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3358____DOLLAR__203513 =  ( n3357____DOLLAR__203510 ) == ( 16'd13 )  ;
assign n3359____DOLLAR__203506 = aes_key[111:104] ;
assign n3360____DOLLAR__203515 =  ( n3358____DOLLAR__203513 ) ? ( ACC ) : ( n3359____DOLLAR__203506 ) ;
assign n3361____DOLLAR__203494 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3362____DOLLAR__203497 =  ( n3361____DOLLAR__203494 ) == ( 16'd12 )  ;
assign n3363____DOLLAR__203490 = aes_key[103:96] ;
assign n3364____DOLLAR__203499 =  ( n3362____DOLLAR__203497 ) ? ( ACC ) : ( n3363____DOLLAR__203490 ) ;
assign n3365____DOLLAR__203478 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3366____DOLLAR__203481 =  ( n3365____DOLLAR__203478 ) == ( 16'd11 )  ;
assign n3367____DOLLAR__203474 = aes_key[95:88] ;
assign n3368____DOLLAR__203483 =  ( n3366____DOLLAR__203481 ) ? ( ACC ) : ( n3367____DOLLAR__203474 ) ;
assign n3369____DOLLAR__203462 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3370____DOLLAR__203465 =  ( n3369____DOLLAR__203462 ) == ( 16'd10 )  ;
assign n3371____DOLLAR__203458 = aes_key[87:80] ;
assign n3372____DOLLAR__203467 =  ( n3370____DOLLAR__203465 ) ? ( ACC ) : ( n3371____DOLLAR__203458 ) ;
assign n3373____DOLLAR__203446 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3374____DOLLAR__203449 =  ( n3373____DOLLAR__203446 ) == ( 16'd9 )  ;
assign n3375____DOLLAR__203442 = aes_key[79:72] ;
assign n3376____DOLLAR__203451 =  ( n3374____DOLLAR__203449 ) ? ( ACC ) : ( n3375____DOLLAR__203442 ) ;
assign n3377____DOLLAR__203430 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3378____DOLLAR__203433 =  ( n3377____DOLLAR__203430 ) == ( 16'd8 )  ;
assign n3379____DOLLAR__203426 = aes_key[71:64] ;
assign n3380____DOLLAR__203435 =  ( n3378____DOLLAR__203433 ) ? ( ACC ) : ( n3379____DOLLAR__203426 ) ;
assign n3381____DOLLAR__203414 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3382____DOLLAR__203417 =  ( n3381____DOLLAR__203414 ) == ( 16'd7 )  ;
assign n3383____DOLLAR__203410 = aes_key[63:56] ;
assign n3384____DOLLAR__203419 =  ( n3382____DOLLAR__203417 ) ? ( ACC ) : ( n3383____DOLLAR__203410 ) ;
assign n3385____DOLLAR__203398 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3386____DOLLAR__203401 =  ( n3385____DOLLAR__203398 ) == ( 16'd6 )  ;
assign n3387____DOLLAR__203394 = aes_key[55:48] ;
assign n3388____DOLLAR__203403 =  ( n3386____DOLLAR__203401 ) ? ( ACC ) : ( n3387____DOLLAR__203394 ) ;
assign n3389____DOLLAR__203382 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3390____DOLLAR__203385 =  ( n3389____DOLLAR__203382 ) == ( 16'd5 )  ;
assign n3391____DOLLAR__203378 = aes_key[47:40] ;
assign n3392____DOLLAR__203387 =  ( n3390____DOLLAR__203385 ) ? ( ACC ) : ( n3391____DOLLAR__203378 ) ;
assign n3393____DOLLAR__203366 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3394____DOLLAR__203369 =  ( n3393____DOLLAR__203366 ) == ( 16'd4 )  ;
assign n3395____DOLLAR__203362 = aes_key[39:32] ;
assign n3396____DOLLAR__203371 =  ( n3394____DOLLAR__203369 ) ? ( ACC ) : ( n3395____DOLLAR__203362 ) ;
assign n3397____DOLLAR__203350 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3398____DOLLAR__203353 =  ( n3397____DOLLAR__203350 ) == ( 16'd3 )  ;
assign n3399____DOLLAR__203346 = aes_key[31:24] ;
assign n3400____DOLLAR__203355 =  ( n3398____DOLLAR__203353 ) ? ( ACC ) : ( n3399____DOLLAR__203346 ) ;
assign n3401____DOLLAR__203334 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3402____DOLLAR__203337 =  ( n3401____DOLLAR__203334 ) == ( 16'd2 )  ;
assign n3403____DOLLAR__203330 = aes_key[23:16] ;
assign n3404____DOLLAR__203339 =  ( n3402____DOLLAR__203337 ) ? ( ACC ) : ( n3403____DOLLAR__203330 ) ;
assign n3405____DOLLAR__203318 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3406____DOLLAR__203321 =  ( n3405____DOLLAR__203318 ) == ( 16'd1 )  ;
assign n3407____DOLLAR__203314 = aes_key[15:8] ;
assign n3408____DOLLAR__203323 =  ( n3406____DOLLAR__203321 ) ? ( ACC ) : ( n3407____DOLLAR__203314 ) ;
assign n3409____DOLLAR__203308 =  ( n3319____DOLLAR__203240 ) - ( 16'd65312 )  ;
assign n3410____DOLLAR__203311 =  ( n3409____DOLLAR__203308 ) == ( 16'd0 )  ;
assign n3411____DOLLAR__203304 = aes_key[7:0] ;
assign n3412____DOLLAR__203313 =  ( n3410____DOLLAR__203311 ) ? ( ACC ) : ( n3411____DOLLAR__203304 ) ;
assign n3413____DOLLAR__203328 =  { ( n3408____DOLLAR__203323 ) , ( n3412____DOLLAR__203313 ) }  ;
assign n3414____DOLLAR__203344 =  { ( n3404____DOLLAR__203339 ) , ( n3413____DOLLAR__203328 ) }  ;
assign n3415____DOLLAR__203360 =  { ( n3400____DOLLAR__203355 ) , ( n3414____DOLLAR__203344 ) }  ;
assign n3416____DOLLAR__203376 =  { ( n3396____DOLLAR__203371 ) , ( n3415____DOLLAR__203360 ) }  ;
assign n3417____DOLLAR__203392 =  { ( n3392____DOLLAR__203387 ) , ( n3416____DOLLAR__203376 ) }  ;
assign n3418____DOLLAR__203408 =  { ( n3388____DOLLAR__203403 ) , ( n3417____DOLLAR__203392 ) }  ;
assign n3419____DOLLAR__203424 =  { ( n3384____DOLLAR__203419 ) , ( n3418____DOLLAR__203408 ) }  ;
assign n3420____DOLLAR__203440 =  { ( n3380____DOLLAR__203435 ) , ( n3419____DOLLAR__203424 ) }  ;
assign n3421____DOLLAR__203456 =  { ( n3376____DOLLAR__203451 ) , ( n3420____DOLLAR__203440 ) }  ;
assign n3422____DOLLAR__203472 =  { ( n3372____DOLLAR__203467 ) , ( n3421____DOLLAR__203456 ) }  ;
assign n3423____DOLLAR__203488 =  { ( n3368____DOLLAR__203483 ) , ( n3422____DOLLAR__203472 ) }  ;
assign n3424____DOLLAR__203504 =  { ( n3364____DOLLAR__203499 ) , ( n3423____DOLLAR__203488 ) }  ;
assign n3425____DOLLAR__203520 =  { ( n3360____DOLLAR__203515 ) , ( n3424____DOLLAR__203504 ) }  ;
assign n3426____DOLLAR__203536 =  { ( n3356____DOLLAR__203531 ) , ( n3425____DOLLAR__203520 ) }  ;
assign n3427____DOLLAR__203552 =  { ( n3352____DOLLAR__203547 ) , ( n3426____DOLLAR__203536 ) }  ;
assign n3428____DOLLAR__203558 =  ( n3348____DOLLAR__203556 ) ? ( n3427____DOLLAR__203552 ) : ( aes_key ) ;
assign n3429____DOLLAR__203811 =  ( aes_status ) == ( 2'd0 )  ;
assign n3430____DOLLAR__203797 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3431____DOLLAR__203800 =  ( n3430____DOLLAR__203797 ) == ( 16'd15 )  ;
assign n3432____DOLLAR__203793 = aes_counter[127:120] ;
assign n3433____DOLLAR__203802 =  ( n3431____DOLLAR__203800 ) ? ( ACC ) : ( n3432____DOLLAR__203793 ) ;
assign n3434____DOLLAR__203781 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3435____DOLLAR__203784 =  ( n3434____DOLLAR__203781 ) == ( 16'd14 )  ;
assign n3436____DOLLAR__203777 = aes_counter[119:112] ;
assign n3437____DOLLAR__203786 =  ( n3435____DOLLAR__203784 ) ? ( ACC ) : ( n3436____DOLLAR__203777 ) ;
assign n3438____DOLLAR__203765 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3439____DOLLAR__203768 =  ( n3438____DOLLAR__203765 ) == ( 16'd13 )  ;
assign n3440____DOLLAR__203761 = aes_counter[111:104] ;
assign n3441____DOLLAR__203770 =  ( n3439____DOLLAR__203768 ) ? ( ACC ) : ( n3440____DOLLAR__203761 ) ;
assign n3442____DOLLAR__203749 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3443____DOLLAR__203752 =  ( n3442____DOLLAR__203749 ) == ( 16'd12 )  ;
assign n3444____DOLLAR__203745 = aes_counter[103:96] ;
assign n3445____DOLLAR__203754 =  ( n3443____DOLLAR__203752 ) ? ( ACC ) : ( n3444____DOLLAR__203745 ) ;
assign n3446____DOLLAR__203733 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3447____DOLLAR__203736 =  ( n3446____DOLLAR__203733 ) == ( 16'd11 )  ;
assign n3448____DOLLAR__203729 = aes_counter[95:88] ;
assign n3449____DOLLAR__203738 =  ( n3447____DOLLAR__203736 ) ? ( ACC ) : ( n3448____DOLLAR__203729 ) ;
assign n3450____DOLLAR__203717 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3451____DOLLAR__203720 =  ( n3450____DOLLAR__203717 ) == ( 16'd10 )  ;
assign n3452____DOLLAR__203713 = aes_counter[87:80] ;
assign n3453____DOLLAR__203722 =  ( n3451____DOLLAR__203720 ) ? ( ACC ) : ( n3452____DOLLAR__203713 ) ;
assign n3454____DOLLAR__203701 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3455____DOLLAR__203704 =  ( n3454____DOLLAR__203701 ) == ( 16'd9 )  ;
assign n3456____DOLLAR__203697 = aes_counter[79:72] ;
assign n3457____DOLLAR__203706 =  ( n3455____DOLLAR__203704 ) ? ( ACC ) : ( n3456____DOLLAR__203697 ) ;
assign n3458____DOLLAR__203685 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3459____DOLLAR__203688 =  ( n3458____DOLLAR__203685 ) == ( 16'd8 )  ;
assign n3460____DOLLAR__203681 = aes_counter[71:64] ;
assign n3461____DOLLAR__203690 =  ( n3459____DOLLAR__203688 ) ? ( ACC ) : ( n3460____DOLLAR__203681 ) ;
assign n3462____DOLLAR__203669 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3463____DOLLAR__203672 =  ( n3462____DOLLAR__203669 ) == ( 16'd7 )  ;
assign n3464____DOLLAR__203665 = aes_counter[63:56] ;
assign n3465____DOLLAR__203674 =  ( n3463____DOLLAR__203672 ) ? ( ACC ) : ( n3464____DOLLAR__203665 ) ;
assign n3466____DOLLAR__203653 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3467____DOLLAR__203656 =  ( n3466____DOLLAR__203653 ) == ( 16'd6 )  ;
assign n3468____DOLLAR__203649 = aes_counter[55:48] ;
assign n3469____DOLLAR__203658 =  ( n3467____DOLLAR__203656 ) ? ( ACC ) : ( n3468____DOLLAR__203649 ) ;
assign n3470____DOLLAR__203637 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3471____DOLLAR__203640 =  ( n3470____DOLLAR__203637 ) == ( 16'd5 )  ;
assign n3472____DOLLAR__203633 = aes_counter[47:40] ;
assign n3473____DOLLAR__203642 =  ( n3471____DOLLAR__203640 ) ? ( ACC ) : ( n3472____DOLLAR__203633 ) ;
assign n3474____DOLLAR__203621 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3475____DOLLAR__203624 =  ( n3474____DOLLAR__203621 ) == ( 16'd4 )  ;
assign n3476____DOLLAR__203617 = aes_counter[39:32] ;
assign n3477____DOLLAR__203626 =  ( n3475____DOLLAR__203624 ) ? ( ACC ) : ( n3476____DOLLAR__203617 ) ;
assign n3478____DOLLAR__203605 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3479____DOLLAR__203608 =  ( n3478____DOLLAR__203605 ) == ( 16'd3 )  ;
assign n3480____DOLLAR__203601 = aes_counter[31:24] ;
assign n3481____DOLLAR__203610 =  ( n3479____DOLLAR__203608 ) ? ( ACC ) : ( n3480____DOLLAR__203601 ) ;
assign n3482____DOLLAR__203589 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3483____DOLLAR__203592 =  ( n3482____DOLLAR__203589 ) == ( 16'd2 )  ;
assign n3484____DOLLAR__203585 = aes_counter[23:16] ;
assign n3485____DOLLAR__203594 =  ( n3483____DOLLAR__203592 ) ? ( ACC ) : ( n3484____DOLLAR__203585 ) ;
assign n3486____DOLLAR__203573 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3487____DOLLAR__203576 =  ( n3486____DOLLAR__203573 ) == ( 16'd1 )  ;
assign n3488____DOLLAR__203569 = aes_counter[15:8] ;
assign n3489____DOLLAR__203578 =  ( n3487____DOLLAR__203576 ) ? ( ACC ) : ( n3488____DOLLAR__203569 ) ;
assign n3490____DOLLAR__203563 =  ( n3319____DOLLAR__203240 ) - ( 16'd65296 )  ;
assign n3491____DOLLAR__203566 =  ( n3490____DOLLAR__203563 ) == ( 16'd0 )  ;
assign n3492____DOLLAR__203559 = aes_counter[7:0] ;
assign n3493____DOLLAR__203568 =  ( n3491____DOLLAR__203566 ) ? ( ACC ) : ( n3492____DOLLAR__203559 ) ;
assign n3494____DOLLAR__203583 =  { ( n3489____DOLLAR__203578 ) , ( n3493____DOLLAR__203568 ) }  ;
assign n3495____DOLLAR__203599 =  { ( n3485____DOLLAR__203594 ) , ( n3494____DOLLAR__203583 ) }  ;
assign n3496____DOLLAR__203615 =  { ( n3481____DOLLAR__203610 ) , ( n3495____DOLLAR__203599 ) }  ;
assign n3497____DOLLAR__203631 =  { ( n3477____DOLLAR__203626 ) , ( n3496____DOLLAR__203615 ) }  ;
assign n3498____DOLLAR__203647 =  { ( n3473____DOLLAR__203642 ) , ( n3497____DOLLAR__203631 ) }  ;
assign n3499____DOLLAR__203663 =  { ( n3469____DOLLAR__203658 ) , ( n3498____DOLLAR__203647 ) }  ;
assign n3500____DOLLAR__203679 =  { ( n3465____DOLLAR__203674 ) , ( n3499____DOLLAR__203663 ) }  ;
assign n3501____DOLLAR__203695 =  { ( n3461____DOLLAR__203690 ) , ( n3500____DOLLAR__203679 ) }  ;
assign n3502____DOLLAR__203711 =  { ( n3457____DOLLAR__203706 ) , ( n3501____DOLLAR__203695 ) }  ;
assign n3503____DOLLAR__203727 =  { ( n3453____DOLLAR__203722 ) , ( n3502____DOLLAR__203711 ) }  ;
assign n3504____DOLLAR__203743 =  { ( n3449____DOLLAR__203738 ) , ( n3503____DOLLAR__203727 ) }  ;
assign n3505____DOLLAR__203759 =  { ( n3445____DOLLAR__203754 ) , ( n3504____DOLLAR__203743 ) }  ;
assign n3506____DOLLAR__203775 =  { ( n3441____DOLLAR__203770 ) , ( n3505____DOLLAR__203759 ) }  ;
assign n3507____DOLLAR__203791 =  { ( n3437____DOLLAR__203786 ) , ( n3506____DOLLAR__203775 ) }  ;
assign n3508____DOLLAR__203807 =  { ( n3433____DOLLAR__203802 ) , ( n3507____DOLLAR__203791 ) }  ;
assign n3509____DOLLAR__203813 =  ( n3429____DOLLAR__203811 ) ? ( n3508____DOLLAR__203807 ) : ( aes_counter ) ;
assign n3510____DOLLAR__203823 =  ( aes_status ) == ( 2'd0 )  ;
assign n3511____DOLLAR__203818 =  ( n3319____DOLLAR__203240 ) == ( 16'd65280 )  ;
assign n3512____DOLLAR__203820 =  ( n3511____DOLLAR__203818 ) ? ( 2'd1 ) : ( aes_status ) ;
assign n3513____DOLLAR__203825 =  ( n3510____DOLLAR__203823 ) ? ( n3512____DOLLAR__203820 ) : ( aes_status ) ;
always @(posedge clk) begin
   if(rst) begin
       ACC <= ACC_randinit ;
       B <= B_randinit ;
       DPH <= DPH_randinit ;
       DPL <= DPL_randinit ;
       IE <= IE_randinit ;
       IP <= IP_randinit ;
       P0 <= P0_randinit ;
       P1 <= P1_randinit ;
       P2 <= P2_randinit ;
       P3 <= P3_randinit ;
       PC <= PC_randinit ;
       PCON <= PCON_randinit ;
       PSW <= PSW_randinit ;
       SBUF <= SBUF_randinit ;
       SCON <= SCON_randinit ;
       SP <= SP_randinit ;
       TCON <= TCON_randinit ;
       TH0 <= TH0_randinit ;
       TH1 <= TH1_randinit ;
       TL0 <= TL0_randinit ;
       TL1 <= TL1_randinit ;
       TMOD <= TMOD_randinit ;
       XRAM_ADDR <= XRAM_ADDR_randinit ;
       XRAM_DATA_IN <= XRAM_DATA_IN_randinit ;
       XRAM_DATA_OUT <= XRAM_DATA_OUT_randinit ;
       oc8051_IRAM_data_0 <= oc8051_IRAM_data_0_randinit ;
       oc8051_IRAM_data_1 <= oc8051_IRAM_data_1_randinit ;
       oc8051_IRAM_data_2 <= oc8051_IRAM_data_2_randinit ;
       oc8051_IRAM_data_3 <= oc8051_IRAM_data_3_randinit ;
       oc8051_IRAM_data_4 <= oc8051_IRAM_data_4_randinit ;
       oc8051_IRAM_data_5 <= oc8051_IRAM_data_5_randinit ;
       oc8051_IRAM_data_6 <= oc8051_IRAM_data_6_randinit ;
       oc8051_IRAM_data_7 <= oc8051_IRAM_data_7_randinit ;
       oc8051_IRAM_data_8 <= oc8051_IRAM_data_8_randinit ;
       oc8051_IRAM_data_9 <= oc8051_IRAM_data_9_randinit ;
       oc8051_IRAM_data_10 <= oc8051_IRAM_data_10_randinit ;
       oc8051_IRAM_data_11 <= oc8051_IRAM_data_11_randinit ;
       oc8051_IRAM_data_12 <= oc8051_IRAM_data_12_randinit ;
       oc8051_IRAM_data_13 <= oc8051_IRAM_data_13_randinit ;
       oc8051_IRAM_data_14 <= oc8051_IRAM_data_14_randinit ;
       oc8051_IRAM_data_15 <= oc8051_IRAM_data_15_randinit ;
       oc8051_ROM_addr_0 <= oc8051_ROM_addr_0_randinit ;
       oc8051_ROM_addr_1 <= oc8051_ROM_addr_1_randinit ;
       oc8051_ROM_addr_2 <= oc8051_ROM_addr_2_randinit ;
       aes_address <= aes_address_randinit ;
       aes_length <= aes_length_randinit ;
       aes_key <= aes_key_randinit ;
       aes_counter <= aes_counter_randinit ;
       aes_status <= aes_status_randinit ;
       __COUNTER_start__n1 <= 0;
   end
   else if(__START__ && __ILA_oc8051_valid__) begin
       if ( __ILA_oc8051_decode_of_I__DOT__240__ ) begin 
           __COUNTER_start__n1 <= 1; end
       else if( (__COUNTER_start__n1 >= 1 ) && ( __COUNTER_start__n1 < 255 )) begin
           __COUNTER_start__n1 <= __COUNTER_start__n1 + 1; end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           ACC <= ACC ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           B <= B ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           DPH <= DPH ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           DPL <= n463____DOLLAR__1232 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           IE <= IE ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           IP <= IP ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           P0 <= P0 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           P1 <= P1 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           P2 <= P2 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           P3 <= n922____DOLLAR__2392 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           PC <= n1513____DOLLAR__3701 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           PCON <= PCON ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           PSW <= PSW ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           SBUF <= SBUF ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           SCON <= SCON ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           SP <= n2213____DOLLAR__5421 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           TCON <= TCON ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           TH0 <= TH0 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           TH1 <= TH1 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           TL0 <= TL0 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           TL1 <= TL1 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           TMOD <= TMOD ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           XRAM_ADDR <= n2800____DOLLAR__6773 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           XRAM_DATA_IN <= XRAM_DATA_IN ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           XRAM_DATA_OUT <= n3312____DOLLAR__8057 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_0 <= oc8051_IRAM_data_0 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_1 <= oc8051_IRAM_data_1 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_2 <= oc8051_IRAM_data_2 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_3 <= oc8051_IRAM_data_3 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_4 <= oc8051_IRAM_data_4 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_5 <= oc8051_IRAM_data_5 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_6 <= oc8051_IRAM_data_6 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_7 <= oc8051_IRAM_data_7 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_8 <= oc8051_IRAM_data_8 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_9 <= oc8051_IRAM_data_9 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_10 <= oc8051_IRAM_data_10 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_11 <= oc8051_IRAM_data_11 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_12 <= oc8051_IRAM_data_12 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_13 <= oc8051_IRAM_data_13 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_14 <= oc8051_IRAM_data_14 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_IRAM_data_15 <= oc8051_IRAM_data_15 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_ROM_addr_0 <= PC ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_ROM_addr_1 <= n3313____DOLLAR__203215 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           oc8051_ROM_addr_2 <= n3314____DOLLAR__203218 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           aes_address <= n3337____DOLLAR__203303 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           aes_length <= n3347____DOLLAR__203272 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           aes_key <= n3428____DOLLAR__203558 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           aes_counter <= n3509____DOLLAR__203813 ;
       end
       if (__ILA_oc8051_decode_of_I__DOT__240__) begin
           aes_status <= n3513____DOLLAR__203825 ;
       end
   end
end
endmodule
