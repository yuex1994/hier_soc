/* PREHEADER */
module fun_sha (
    input [511:0] arg0,
    output [159:0] result
);
//TODO: Add the specific function HERE.
endmodule

/* END OF PREHEADER */
module sha(
__ILA_sha_grant__,
clk,
cmd,
cmdaddr,
cmddata,
rst,
__ILA_sha_acc_decode__,
__ILA_sha_decode_of_I__DOT__0__,
__ILA_sha_decode_of_I__DOT__100__,
__ILA_sha_decode_of_I__DOT__101__,
__ILA_sha_decode_of_I__DOT__102__,
__ILA_sha_decode_of_I__DOT__103__,
__ILA_sha_decode_of_I__DOT__104__,
__ILA_sha_decode_of_I__DOT__105__,
__ILA_sha_decode_of_I__DOT__106__,
__ILA_sha_decode_of_I__DOT__107__,
__ILA_sha_decode_of_I__DOT__108__,
__ILA_sha_decode_of_I__DOT__109__,
__ILA_sha_decode_of_I__DOT__10__,
__ILA_sha_decode_of_I__DOT__110__,
__ILA_sha_decode_of_I__DOT__111__,
__ILA_sha_decode_of_I__DOT__112__,
__ILA_sha_decode_of_I__DOT__113__,
__ILA_sha_decode_of_I__DOT__114__,
__ILA_sha_decode_of_I__DOT__115__,
__ILA_sha_decode_of_I__DOT__116__,
__ILA_sha_decode_of_I__DOT__117__,
__ILA_sha_decode_of_I__DOT__118__,
__ILA_sha_decode_of_I__DOT__119__,
__ILA_sha_decode_of_I__DOT__11__,
__ILA_sha_decode_of_I__DOT__120__,
__ILA_sha_decode_of_I__DOT__121__,
__ILA_sha_decode_of_I__DOT__122__,
__ILA_sha_decode_of_I__DOT__123__,
__ILA_sha_decode_of_I__DOT__124__,
__ILA_sha_decode_of_I__DOT__125__,
__ILA_sha_decode_of_I__DOT__126__,
__ILA_sha_decode_of_I__DOT__127__,
__ILA_sha_decode_of_I__DOT__128__,
__ILA_sha_decode_of_I__DOT__129__,
__ILA_sha_decode_of_I__DOT__12__,
__ILA_sha_decode_of_I__DOT__130__,
__ILA_sha_decode_of_I__DOT__131__,
__ILA_sha_decode_of_I__DOT__132__,
__ILA_sha_decode_of_I__DOT__133__,
__ILA_sha_decode_of_I__DOT__134__,
__ILA_sha_decode_of_I__DOT__135__,
__ILA_sha_decode_of_I__DOT__136__,
__ILA_sha_decode_of_I__DOT__137__,
__ILA_sha_decode_of_I__DOT__138__,
__ILA_sha_decode_of_I__DOT__139__,
__ILA_sha_decode_of_I__DOT__13__,
__ILA_sha_decode_of_I__DOT__140__,
__ILA_sha_decode_of_I__DOT__141__,
__ILA_sha_decode_of_I__DOT__142__,
__ILA_sha_decode_of_I__DOT__143__,
__ILA_sha_decode_of_I__DOT__144__,
__ILA_sha_decode_of_I__DOT__145__,
__ILA_sha_decode_of_I__DOT__146__,
__ILA_sha_decode_of_I__DOT__147__,
__ILA_sha_decode_of_I__DOT__148__,
__ILA_sha_decode_of_I__DOT__149__,
__ILA_sha_decode_of_I__DOT__14__,
__ILA_sha_decode_of_I__DOT__150__,
__ILA_sha_decode_of_I__DOT__151__,
__ILA_sha_decode_of_I__DOT__152__,
__ILA_sha_decode_of_I__DOT__153__,
__ILA_sha_decode_of_I__DOT__154__,
__ILA_sha_decode_of_I__DOT__155__,
__ILA_sha_decode_of_I__DOT__156__,
__ILA_sha_decode_of_I__DOT__157__,
__ILA_sha_decode_of_I__DOT__158__,
__ILA_sha_decode_of_I__DOT__159__,
__ILA_sha_decode_of_I__DOT__15__,
__ILA_sha_decode_of_I__DOT__16__,
__ILA_sha_decode_of_I__DOT__17__,
__ILA_sha_decode_of_I__DOT__18__,
__ILA_sha_decode_of_I__DOT__19__,
__ILA_sha_decode_of_I__DOT__1__,
__ILA_sha_decode_of_I__DOT__20__,
__ILA_sha_decode_of_I__DOT__21__,
__ILA_sha_decode_of_I__DOT__22__,
__ILA_sha_decode_of_I__DOT__23__,
__ILA_sha_decode_of_I__DOT__24__,
__ILA_sha_decode_of_I__DOT__25__,
__ILA_sha_decode_of_I__DOT__26__,
__ILA_sha_decode_of_I__DOT__27__,
__ILA_sha_decode_of_I__DOT__28__,
__ILA_sha_decode_of_I__DOT__29__,
__ILA_sha_decode_of_I__DOT__2__,
__ILA_sha_decode_of_I__DOT__30__,
__ILA_sha_decode_of_I__DOT__31__,
__ILA_sha_decode_of_I__DOT__32__,
__ILA_sha_decode_of_I__DOT__33__,
__ILA_sha_decode_of_I__DOT__34__,
__ILA_sha_decode_of_I__DOT__35__,
__ILA_sha_decode_of_I__DOT__36__,
__ILA_sha_decode_of_I__DOT__37__,
__ILA_sha_decode_of_I__DOT__38__,
__ILA_sha_decode_of_I__DOT__39__,
__ILA_sha_decode_of_I__DOT__3__,
__ILA_sha_decode_of_I__DOT__40__,
__ILA_sha_decode_of_I__DOT__41__,
__ILA_sha_decode_of_I__DOT__42__,
__ILA_sha_decode_of_I__DOT__43__,
__ILA_sha_decode_of_I__DOT__44__,
__ILA_sha_decode_of_I__DOT__45__,
__ILA_sha_decode_of_I__DOT__46__,
__ILA_sha_decode_of_I__DOT__47__,
__ILA_sha_decode_of_I__DOT__48__,
__ILA_sha_decode_of_I__DOT__49__,
__ILA_sha_decode_of_I__DOT__4__,
__ILA_sha_decode_of_I__DOT__50__,
__ILA_sha_decode_of_I__DOT__51__,
__ILA_sha_decode_of_I__DOT__52__,
__ILA_sha_decode_of_I__DOT__53__,
__ILA_sha_decode_of_I__DOT__54__,
__ILA_sha_decode_of_I__DOT__55__,
__ILA_sha_decode_of_I__DOT__56__,
__ILA_sha_decode_of_I__DOT__57__,
__ILA_sha_decode_of_I__DOT__58__,
__ILA_sha_decode_of_I__DOT__59__,
__ILA_sha_decode_of_I__DOT__5__,
__ILA_sha_decode_of_I__DOT__60__,
__ILA_sha_decode_of_I__DOT__61__,
__ILA_sha_decode_of_I__DOT__62__,
__ILA_sha_decode_of_I__DOT__63__,
__ILA_sha_decode_of_I__DOT__64__,
__ILA_sha_decode_of_I__DOT__65__,
__ILA_sha_decode_of_I__DOT__66__,
__ILA_sha_decode_of_I__DOT__67__,
__ILA_sha_decode_of_I__DOT__68__,
__ILA_sha_decode_of_I__DOT__69__,
__ILA_sha_decode_of_I__DOT__6__,
__ILA_sha_decode_of_I__DOT__70__,
__ILA_sha_decode_of_I__DOT__71__,
__ILA_sha_decode_of_I__DOT__72__,
__ILA_sha_decode_of_I__DOT__73__,
__ILA_sha_decode_of_I__DOT__74__,
__ILA_sha_decode_of_I__DOT__75__,
__ILA_sha_decode_of_I__DOT__76__,
__ILA_sha_decode_of_I__DOT__77__,
__ILA_sha_decode_of_I__DOT__78__,
__ILA_sha_decode_of_I__DOT__79__,
__ILA_sha_decode_of_I__DOT__7__,
__ILA_sha_decode_of_I__DOT__80__,
__ILA_sha_decode_of_I__DOT__81__,
__ILA_sha_decode_of_I__DOT__82__,
__ILA_sha_decode_of_I__DOT__83__,
__ILA_sha_decode_of_I__DOT__84__,
__ILA_sha_decode_of_I__DOT__85__,
__ILA_sha_decode_of_I__DOT__86__,
__ILA_sha_decode_of_I__DOT__87__,
__ILA_sha_decode_of_I__DOT__88__,
__ILA_sha_decode_of_I__DOT__89__,
__ILA_sha_decode_of_I__DOT__8__,
__ILA_sha_decode_of_I__DOT__90__,
__ILA_sha_decode_of_I__DOT__91__,
__ILA_sha_decode_of_I__DOT__92__,
__ILA_sha_decode_of_I__DOT__93__,
__ILA_sha_decode_of_I__DOT__94__,
__ILA_sha_decode_of_I__DOT__95__,
__ILA_sha_decode_of_I__DOT__96__,
__ILA_sha_decode_of_I__DOT__97__,
__ILA_sha_decode_of_I__DOT__98__,
__ILA_sha_decode_of_I__DOT__99__,
__ILA_sha_decode_of_I__DOT__9__,
__ILA_sha_valid__,
XRAM_data_n915,
XRAM_data_n919,
XRAM_data_n924,
XRAM_data_n929,
XRAM_data_n934,
XRAM_data_n939,
XRAM_data_n944,
XRAM_data_n949,
XRAM_data_n954,
XRAM_data_n959,
XRAM_data_n964,
XRAM_data_n969,
XRAM_data_n974,
XRAM_data_n979,
XRAM_data_n984,
XRAM_data_n989,
XRAM_data_n994,
XRAM_data_n999,
XRAM_data_n1004,
XRAM_data_n1009,
XRAM_data_n1014,
XRAM_data_n1019,
XRAM_data_n1024,
XRAM_data_n1029,
XRAM_data_n1034,
XRAM_data_n1039,
XRAM_data_n1044,
XRAM_data_n1049,
XRAM_data_n1054,
XRAM_data_n1059,
XRAM_data_n1064,
XRAM_data_n1069,
XRAM_data_n1074,
XRAM_data_n1079,
XRAM_data_n1084,
XRAM_data_n1089,
XRAM_data_n1094,
XRAM_data_n1099,
XRAM_data_n1104,
XRAM_data_n1109,
XRAM_data_n1114,
XRAM_data_n1119,
XRAM_data_n1124,
XRAM_data_n1129,
XRAM_data_n1134,
XRAM_data_n1139,
XRAM_data_n1144,
XRAM_data_n1149,
XRAM_data_n1154,
XRAM_data_n1159,
XRAM_data_n1164,
XRAM_data_n1169,
XRAM_data_n1174,
XRAM_data_n1179,
XRAM_data_n1184,
XRAM_data_n1189,
XRAM_data_n1194,
XRAM_data_n1199,
XRAM_data_n1204,
XRAM_data_n1209,
XRAM_data_n1214,
XRAM_data_n1219,
XRAM_data_n1224,
XRAM_data_n1229,
XRAM_addr_n914,
XRAM_addr_n918,
XRAM_addr_n923,
XRAM_addr_n928,
XRAM_addr_n933,
XRAM_addr_n938,
XRAM_addr_n943,
XRAM_addr_n948,
XRAM_addr_n953,
XRAM_addr_n958,
XRAM_addr_n963,
XRAM_addr_n968,
XRAM_addr_n973,
XRAM_addr_n978,
XRAM_addr_n983,
XRAM_addr_n988,
XRAM_addr_n993,
XRAM_addr_n998,
XRAM_addr_n1003,
XRAM_addr_n1008,
XRAM_addr_n1013,
XRAM_addr_n1018,
XRAM_addr_n1023,
XRAM_addr_n1028,
XRAM_addr_n1033,
XRAM_addr_n1038,
XRAM_addr_n1043,
XRAM_addr_n1048,
XRAM_addr_n1053,
XRAM_addr_n1058,
XRAM_addr_n1063,
XRAM_addr_n1068,
XRAM_addr_n1073,
XRAM_addr_n1078,
XRAM_addr_n1083,
XRAM_addr_n1088,
XRAM_addr_n1093,
XRAM_addr_n1098,
XRAM_addr_n1103,
XRAM_addr_n1108,
XRAM_addr_n1113,
XRAM_addr_n1118,
XRAM_addr_n1123,
XRAM_addr_n1128,
XRAM_addr_n1133,
XRAM_addr_n1138,
XRAM_addr_n1143,
XRAM_addr_n1148,
XRAM_addr_n1153,
XRAM_addr_n1158,
XRAM_addr_n1163,
XRAM_addr_n1168,
XRAM_addr_n1173,
XRAM_addr_n1178,
XRAM_addr_n1183,
XRAM_addr_n1188,
XRAM_addr_n1193,
XRAM_addr_n1198,
XRAM_addr_n1203,
XRAM_addr_n1208,
XRAM_addr_n1213,
XRAM_addr_n1218,
XRAM_addr_n1223,
XRAM_addr_n1228,
XRAM_addr0,
XRAM_data0,
XRAM_wen0,
XRAM_addr1,
XRAM_data1,
XRAM_wen1,
XRAM_addr2,
XRAM_data2,
XRAM_wen2,
XRAM_addr3,
XRAM_data3,
XRAM_wen3,
XRAM_addr4,
XRAM_data4,
XRAM_wen4,
XRAM_addr5,
XRAM_data5,
XRAM_wen5,
XRAM_addr6,
XRAM_data6,
XRAM_wen6,
XRAM_addr7,
XRAM_data7,
XRAM_wen7,
dataout,
sha_bytes_read,
sha_hs_data,
sha_len,
sha_rd_data,
sha_rdaddr,
sha_state,
sha_wraddr
);
input    [159:0] __ILA_sha_grant__;
input            clk;
input      [1:0] cmd;
input     [15:0] cmdaddr;
input      [7:0] cmddata;
input            rst;
input      [7:0] XRAM_data_n915;
input      [7:0] XRAM_data_n919;
input      [7:0] XRAM_data_n924;
input      [7:0] XRAM_data_n929;
input      [7:0] XRAM_data_n934;
input      [7:0] XRAM_data_n939;
input      [7:0] XRAM_data_n944;
input      [7:0] XRAM_data_n949;
input      [7:0] XRAM_data_n954;
input      [7:0] XRAM_data_n959;
input      [7:0] XRAM_data_n964;
input      [7:0] XRAM_data_n969;
input      [7:0] XRAM_data_n974;
input      [7:0] XRAM_data_n979;
input      [7:0] XRAM_data_n984;
input      [7:0] XRAM_data_n989;
input      [7:0] XRAM_data_n994;
input      [7:0] XRAM_data_n999;
input      [7:0] XRAM_data_n1004;
input      [7:0] XRAM_data_n1009;
input      [7:0] XRAM_data_n1014;
input      [7:0] XRAM_data_n1019;
input      [7:0] XRAM_data_n1024;
input      [7:0] XRAM_data_n1029;
input      [7:0] XRAM_data_n1034;
input      [7:0] XRAM_data_n1039;
input      [7:0] XRAM_data_n1044;
input      [7:0] XRAM_data_n1049;
input      [7:0] XRAM_data_n1054;
input      [7:0] XRAM_data_n1059;
input      [7:0] XRAM_data_n1064;
input      [7:0] XRAM_data_n1069;
input      [7:0] XRAM_data_n1074;
input      [7:0] XRAM_data_n1079;
input      [7:0] XRAM_data_n1084;
input      [7:0] XRAM_data_n1089;
input      [7:0] XRAM_data_n1094;
input      [7:0] XRAM_data_n1099;
input      [7:0] XRAM_data_n1104;
input      [7:0] XRAM_data_n1109;
input      [7:0] XRAM_data_n1114;
input      [7:0] XRAM_data_n1119;
input      [7:0] XRAM_data_n1124;
input      [7:0] XRAM_data_n1129;
input      [7:0] XRAM_data_n1134;
input      [7:0] XRAM_data_n1139;
input      [7:0] XRAM_data_n1144;
input      [7:0] XRAM_data_n1149;
input      [7:0] XRAM_data_n1154;
input      [7:0] XRAM_data_n1159;
input      [7:0] XRAM_data_n1164;
input      [7:0] XRAM_data_n1169;
input      [7:0] XRAM_data_n1174;
input      [7:0] XRAM_data_n1179;
input      [7:0] XRAM_data_n1184;
input      [7:0] XRAM_data_n1189;
input      [7:0] XRAM_data_n1194;
input      [7:0] XRAM_data_n1199;
input      [7:0] XRAM_data_n1204;
input      [7:0] XRAM_data_n1209;
input      [7:0] XRAM_data_n1214;
input      [7:0] XRAM_data_n1219;
input      [7:0] XRAM_data_n1224;
input      [7:0] XRAM_data_n1229;
output    [159:0] __ILA_sha_acc_decode__;
output            __ILA_sha_decode_of_I__DOT__0__;
output            __ILA_sha_decode_of_I__DOT__100__;
output            __ILA_sha_decode_of_I__DOT__101__;
output            __ILA_sha_decode_of_I__DOT__102__;
output            __ILA_sha_decode_of_I__DOT__103__;
output            __ILA_sha_decode_of_I__DOT__104__;
output            __ILA_sha_decode_of_I__DOT__105__;
output            __ILA_sha_decode_of_I__DOT__106__;
output            __ILA_sha_decode_of_I__DOT__107__;
output            __ILA_sha_decode_of_I__DOT__108__;
output            __ILA_sha_decode_of_I__DOT__109__;
output            __ILA_sha_decode_of_I__DOT__10__;
output            __ILA_sha_decode_of_I__DOT__110__;
output            __ILA_sha_decode_of_I__DOT__111__;
output            __ILA_sha_decode_of_I__DOT__112__;
output            __ILA_sha_decode_of_I__DOT__113__;
output            __ILA_sha_decode_of_I__DOT__114__;
output            __ILA_sha_decode_of_I__DOT__115__;
output            __ILA_sha_decode_of_I__DOT__116__;
output            __ILA_sha_decode_of_I__DOT__117__;
output            __ILA_sha_decode_of_I__DOT__118__;
output            __ILA_sha_decode_of_I__DOT__119__;
output            __ILA_sha_decode_of_I__DOT__11__;
output            __ILA_sha_decode_of_I__DOT__120__;
output            __ILA_sha_decode_of_I__DOT__121__;
output            __ILA_sha_decode_of_I__DOT__122__;
output            __ILA_sha_decode_of_I__DOT__123__;
output            __ILA_sha_decode_of_I__DOT__124__;
output            __ILA_sha_decode_of_I__DOT__125__;
output            __ILA_sha_decode_of_I__DOT__126__;
output            __ILA_sha_decode_of_I__DOT__127__;
output            __ILA_sha_decode_of_I__DOT__128__;
output            __ILA_sha_decode_of_I__DOT__129__;
output            __ILA_sha_decode_of_I__DOT__12__;
output            __ILA_sha_decode_of_I__DOT__130__;
output            __ILA_sha_decode_of_I__DOT__131__;
output            __ILA_sha_decode_of_I__DOT__132__;
output            __ILA_sha_decode_of_I__DOT__133__;
output            __ILA_sha_decode_of_I__DOT__134__;
output            __ILA_sha_decode_of_I__DOT__135__;
output            __ILA_sha_decode_of_I__DOT__136__;
output            __ILA_sha_decode_of_I__DOT__137__;
output            __ILA_sha_decode_of_I__DOT__138__;
output            __ILA_sha_decode_of_I__DOT__139__;
output            __ILA_sha_decode_of_I__DOT__13__;
output            __ILA_sha_decode_of_I__DOT__140__;
output            __ILA_sha_decode_of_I__DOT__141__;
output            __ILA_sha_decode_of_I__DOT__142__;
output            __ILA_sha_decode_of_I__DOT__143__;
output            __ILA_sha_decode_of_I__DOT__144__;
output            __ILA_sha_decode_of_I__DOT__145__;
output            __ILA_sha_decode_of_I__DOT__146__;
output            __ILA_sha_decode_of_I__DOT__147__;
output            __ILA_sha_decode_of_I__DOT__148__;
output            __ILA_sha_decode_of_I__DOT__149__;
output            __ILA_sha_decode_of_I__DOT__14__;
output            __ILA_sha_decode_of_I__DOT__150__;
output            __ILA_sha_decode_of_I__DOT__151__;
output            __ILA_sha_decode_of_I__DOT__152__;
output            __ILA_sha_decode_of_I__DOT__153__;
output            __ILA_sha_decode_of_I__DOT__154__;
output            __ILA_sha_decode_of_I__DOT__155__;
output            __ILA_sha_decode_of_I__DOT__156__;
output            __ILA_sha_decode_of_I__DOT__157__;
output            __ILA_sha_decode_of_I__DOT__158__;
output            __ILA_sha_decode_of_I__DOT__159__;
output            __ILA_sha_decode_of_I__DOT__15__;
output            __ILA_sha_decode_of_I__DOT__16__;
output            __ILA_sha_decode_of_I__DOT__17__;
output            __ILA_sha_decode_of_I__DOT__18__;
output            __ILA_sha_decode_of_I__DOT__19__;
output            __ILA_sha_decode_of_I__DOT__1__;
output            __ILA_sha_decode_of_I__DOT__20__;
output            __ILA_sha_decode_of_I__DOT__21__;
output            __ILA_sha_decode_of_I__DOT__22__;
output            __ILA_sha_decode_of_I__DOT__23__;
output            __ILA_sha_decode_of_I__DOT__24__;
output            __ILA_sha_decode_of_I__DOT__25__;
output            __ILA_sha_decode_of_I__DOT__26__;
output            __ILA_sha_decode_of_I__DOT__27__;
output            __ILA_sha_decode_of_I__DOT__28__;
output            __ILA_sha_decode_of_I__DOT__29__;
output            __ILA_sha_decode_of_I__DOT__2__;
output            __ILA_sha_decode_of_I__DOT__30__;
output            __ILA_sha_decode_of_I__DOT__31__;
output            __ILA_sha_decode_of_I__DOT__32__;
output            __ILA_sha_decode_of_I__DOT__33__;
output            __ILA_sha_decode_of_I__DOT__34__;
output            __ILA_sha_decode_of_I__DOT__35__;
output            __ILA_sha_decode_of_I__DOT__36__;
output            __ILA_sha_decode_of_I__DOT__37__;
output            __ILA_sha_decode_of_I__DOT__38__;
output            __ILA_sha_decode_of_I__DOT__39__;
output            __ILA_sha_decode_of_I__DOT__3__;
output            __ILA_sha_decode_of_I__DOT__40__;
output            __ILA_sha_decode_of_I__DOT__41__;
output            __ILA_sha_decode_of_I__DOT__42__;
output            __ILA_sha_decode_of_I__DOT__43__;
output            __ILA_sha_decode_of_I__DOT__44__;
output            __ILA_sha_decode_of_I__DOT__45__;
output            __ILA_sha_decode_of_I__DOT__46__;
output            __ILA_sha_decode_of_I__DOT__47__;
output            __ILA_sha_decode_of_I__DOT__48__;
output            __ILA_sha_decode_of_I__DOT__49__;
output            __ILA_sha_decode_of_I__DOT__4__;
output            __ILA_sha_decode_of_I__DOT__50__;
output            __ILA_sha_decode_of_I__DOT__51__;
output            __ILA_sha_decode_of_I__DOT__52__;
output            __ILA_sha_decode_of_I__DOT__53__;
output            __ILA_sha_decode_of_I__DOT__54__;
output            __ILA_sha_decode_of_I__DOT__55__;
output            __ILA_sha_decode_of_I__DOT__56__;
output            __ILA_sha_decode_of_I__DOT__57__;
output            __ILA_sha_decode_of_I__DOT__58__;
output            __ILA_sha_decode_of_I__DOT__59__;
output            __ILA_sha_decode_of_I__DOT__5__;
output            __ILA_sha_decode_of_I__DOT__60__;
output            __ILA_sha_decode_of_I__DOT__61__;
output            __ILA_sha_decode_of_I__DOT__62__;
output            __ILA_sha_decode_of_I__DOT__63__;
output            __ILA_sha_decode_of_I__DOT__64__;
output            __ILA_sha_decode_of_I__DOT__65__;
output            __ILA_sha_decode_of_I__DOT__66__;
output            __ILA_sha_decode_of_I__DOT__67__;
output            __ILA_sha_decode_of_I__DOT__68__;
output            __ILA_sha_decode_of_I__DOT__69__;
output            __ILA_sha_decode_of_I__DOT__6__;
output            __ILA_sha_decode_of_I__DOT__70__;
output            __ILA_sha_decode_of_I__DOT__71__;
output            __ILA_sha_decode_of_I__DOT__72__;
output            __ILA_sha_decode_of_I__DOT__73__;
output            __ILA_sha_decode_of_I__DOT__74__;
output            __ILA_sha_decode_of_I__DOT__75__;
output            __ILA_sha_decode_of_I__DOT__76__;
output            __ILA_sha_decode_of_I__DOT__77__;
output            __ILA_sha_decode_of_I__DOT__78__;
output            __ILA_sha_decode_of_I__DOT__79__;
output            __ILA_sha_decode_of_I__DOT__7__;
output            __ILA_sha_decode_of_I__DOT__80__;
output            __ILA_sha_decode_of_I__DOT__81__;
output            __ILA_sha_decode_of_I__DOT__82__;
output            __ILA_sha_decode_of_I__DOT__83__;
output            __ILA_sha_decode_of_I__DOT__84__;
output            __ILA_sha_decode_of_I__DOT__85__;
output            __ILA_sha_decode_of_I__DOT__86__;
output            __ILA_sha_decode_of_I__DOT__87__;
output            __ILA_sha_decode_of_I__DOT__88__;
output            __ILA_sha_decode_of_I__DOT__89__;
output            __ILA_sha_decode_of_I__DOT__8__;
output            __ILA_sha_decode_of_I__DOT__90__;
output            __ILA_sha_decode_of_I__DOT__91__;
output            __ILA_sha_decode_of_I__DOT__92__;
output            __ILA_sha_decode_of_I__DOT__93__;
output            __ILA_sha_decode_of_I__DOT__94__;
output            __ILA_sha_decode_of_I__DOT__95__;
output            __ILA_sha_decode_of_I__DOT__96__;
output            __ILA_sha_decode_of_I__DOT__97__;
output            __ILA_sha_decode_of_I__DOT__98__;
output            __ILA_sha_decode_of_I__DOT__99__;
output            __ILA_sha_decode_of_I__DOT__9__;
output            __ILA_sha_valid__;
output     [15:0] XRAM_addr_n914;
output     [15:0] XRAM_addr_n918;
output     [15:0] XRAM_addr_n923;
output     [15:0] XRAM_addr_n928;
output     [15:0] XRAM_addr_n933;
output     [15:0] XRAM_addr_n938;
output     [15:0] XRAM_addr_n943;
output     [15:0] XRAM_addr_n948;
output     [15:0] XRAM_addr_n953;
output     [15:0] XRAM_addr_n958;
output     [15:0] XRAM_addr_n963;
output     [15:0] XRAM_addr_n968;
output     [15:0] XRAM_addr_n973;
output     [15:0] XRAM_addr_n978;
output     [15:0] XRAM_addr_n983;
output     [15:0] XRAM_addr_n988;
output     [15:0] XRAM_addr_n993;
output     [15:0] XRAM_addr_n998;
output     [15:0] XRAM_addr_n1003;
output     [15:0] XRAM_addr_n1008;
output     [15:0] XRAM_addr_n1013;
output     [15:0] XRAM_addr_n1018;
output     [15:0] XRAM_addr_n1023;
output     [15:0] XRAM_addr_n1028;
output     [15:0] XRAM_addr_n1033;
output     [15:0] XRAM_addr_n1038;
output     [15:0] XRAM_addr_n1043;
output     [15:0] XRAM_addr_n1048;
output     [15:0] XRAM_addr_n1053;
output     [15:0] XRAM_addr_n1058;
output     [15:0] XRAM_addr_n1063;
output     [15:0] XRAM_addr_n1068;
output     [15:0] XRAM_addr_n1073;
output     [15:0] XRAM_addr_n1078;
output     [15:0] XRAM_addr_n1083;
output     [15:0] XRAM_addr_n1088;
output     [15:0] XRAM_addr_n1093;
output     [15:0] XRAM_addr_n1098;
output     [15:0] XRAM_addr_n1103;
output     [15:0] XRAM_addr_n1108;
output     [15:0] XRAM_addr_n1113;
output     [15:0] XRAM_addr_n1118;
output     [15:0] XRAM_addr_n1123;
output     [15:0] XRAM_addr_n1128;
output     [15:0] XRAM_addr_n1133;
output     [15:0] XRAM_addr_n1138;
output     [15:0] XRAM_addr_n1143;
output     [15:0] XRAM_addr_n1148;
output     [15:0] XRAM_addr_n1153;
output     [15:0] XRAM_addr_n1158;
output     [15:0] XRAM_addr_n1163;
output     [15:0] XRAM_addr_n1168;
output     [15:0] XRAM_addr_n1173;
output     [15:0] XRAM_addr_n1178;
output     [15:0] XRAM_addr_n1183;
output     [15:0] XRAM_addr_n1188;
output     [15:0] XRAM_addr_n1193;
output     [15:0] XRAM_addr_n1198;
output     [15:0] XRAM_addr_n1203;
output     [15:0] XRAM_addr_n1208;
output     [15:0] XRAM_addr_n1213;
output     [15:0] XRAM_addr_n1218;
output     [15:0] XRAM_addr_n1223;
output     [15:0] XRAM_addr_n1228;
output     [15:0] XRAM_addr0;
output      [7:0] XRAM_data0;
output            XRAM_wen0;
output     [15:0] XRAM_addr1;
output      [7:0] XRAM_data1;
output            XRAM_wen1;
output     [15:0] XRAM_addr2;
output      [7:0] XRAM_data2;
output            XRAM_wen2;
output     [15:0] XRAM_addr3;
output      [7:0] XRAM_data3;
output            XRAM_wen3;
output     [15:0] XRAM_addr4;
output      [7:0] XRAM_data4;
output            XRAM_wen4;
output     [15:0] XRAM_addr5;
output      [7:0] XRAM_data5;
output            XRAM_wen5;
output     [15:0] XRAM_addr6;
output      [7:0] XRAM_data6;
output            XRAM_wen6;
output     [15:0] XRAM_addr7;
output      [7:0] XRAM_data7;
output            XRAM_wen7;
output reg      [7:0] dataout;
output reg     [15:0] sha_bytes_read;
output reg    [159:0] sha_hs_data;
output reg     [15:0] sha_len;
output reg    [511:0] sha_rd_data;
output reg     [15:0] sha_rdaddr;
output reg      [2:0] sha_state;
output reg     [15:0] sha_wraddr;
wire     [15:0] XRAM_addr0;
wire     [15:0] XRAM_addr1;
wire     [15:0] XRAM_addr2;
wire     [15:0] XRAM_addr3;
wire     [15:0] XRAM_addr4;
wire     [15:0] XRAM_addr5;
wire     [15:0] XRAM_addr6;
wire     [15:0] XRAM_addr7;
wire     [15:0] XRAM_addr_n1003;
wire     [15:0] XRAM_addr_n1008;
wire     [15:0] XRAM_addr_n1013;
wire     [15:0] XRAM_addr_n1018;
wire     [15:0] XRAM_addr_n1023;
wire     [15:0] XRAM_addr_n1028;
wire     [15:0] XRAM_addr_n1033;
wire     [15:0] XRAM_addr_n1038;
wire     [15:0] XRAM_addr_n1043;
wire     [15:0] XRAM_addr_n1048;
wire     [15:0] XRAM_addr_n1053;
wire     [15:0] XRAM_addr_n1058;
wire     [15:0] XRAM_addr_n1063;
wire     [15:0] XRAM_addr_n1068;
wire     [15:0] XRAM_addr_n1073;
wire     [15:0] XRAM_addr_n1078;
wire     [15:0] XRAM_addr_n1083;
wire     [15:0] XRAM_addr_n1088;
wire     [15:0] XRAM_addr_n1093;
wire     [15:0] XRAM_addr_n1098;
wire     [15:0] XRAM_addr_n1103;
wire     [15:0] XRAM_addr_n1108;
wire     [15:0] XRAM_addr_n1113;
wire     [15:0] XRAM_addr_n1118;
wire     [15:0] XRAM_addr_n1123;
wire     [15:0] XRAM_addr_n1128;
wire     [15:0] XRAM_addr_n1133;
wire     [15:0] XRAM_addr_n1138;
wire     [15:0] XRAM_addr_n1143;
wire     [15:0] XRAM_addr_n1148;
wire     [15:0] XRAM_addr_n1153;
wire     [15:0] XRAM_addr_n1158;
wire     [15:0] XRAM_addr_n1163;
wire     [15:0] XRAM_addr_n1168;
wire     [15:0] XRAM_addr_n1173;
wire     [15:0] XRAM_addr_n1178;
wire     [15:0] XRAM_addr_n1183;
wire     [15:0] XRAM_addr_n1188;
wire     [15:0] XRAM_addr_n1193;
wire     [15:0] XRAM_addr_n1198;
wire     [15:0] XRAM_addr_n1203;
wire     [15:0] XRAM_addr_n1208;
wire     [15:0] XRAM_addr_n1213;
wire     [15:0] XRAM_addr_n1218;
wire     [15:0] XRAM_addr_n1223;
wire     [15:0] XRAM_addr_n1228;
wire     [15:0] XRAM_addr_n914;
wire     [15:0] XRAM_addr_n918;
wire     [15:0] XRAM_addr_n923;
wire     [15:0] XRAM_addr_n928;
wire     [15:0] XRAM_addr_n933;
wire     [15:0] XRAM_addr_n938;
wire     [15:0] XRAM_addr_n943;
wire     [15:0] XRAM_addr_n948;
wire     [15:0] XRAM_addr_n953;
wire     [15:0] XRAM_addr_n958;
wire     [15:0] XRAM_addr_n963;
wire     [15:0] XRAM_addr_n968;
wire     [15:0] XRAM_addr_n973;
wire     [15:0] XRAM_addr_n978;
wire     [15:0] XRAM_addr_n983;
wire     [15:0] XRAM_addr_n988;
wire     [15:0] XRAM_addr_n993;
wire     [15:0] XRAM_addr_n998;
wire      [7:0] XRAM_data0;
wire      [7:0] XRAM_data1;
wire      [7:0] XRAM_data2;
wire      [7:0] XRAM_data3;
wire      [7:0] XRAM_data4;
wire      [7:0] XRAM_data5;
wire      [7:0] XRAM_data6;
wire      [7:0] XRAM_data7;
wire      [7:0] XRAM_data_n1004;
wire      [7:0] XRAM_data_n1009;
wire      [7:0] XRAM_data_n1014;
wire      [7:0] XRAM_data_n1019;
wire      [7:0] XRAM_data_n1024;
wire      [7:0] XRAM_data_n1029;
wire      [7:0] XRAM_data_n1034;
wire      [7:0] XRAM_data_n1039;
wire      [7:0] XRAM_data_n1044;
wire      [7:0] XRAM_data_n1049;
wire      [7:0] XRAM_data_n1054;
wire      [7:0] XRAM_data_n1059;
wire      [7:0] XRAM_data_n1064;
wire      [7:0] XRAM_data_n1069;
wire      [7:0] XRAM_data_n1074;
wire      [7:0] XRAM_data_n1079;
wire      [7:0] XRAM_data_n1084;
wire      [7:0] XRAM_data_n1089;
wire      [7:0] XRAM_data_n1094;
wire      [7:0] XRAM_data_n1099;
wire      [7:0] XRAM_data_n1104;
wire      [7:0] XRAM_data_n1109;
wire      [7:0] XRAM_data_n1114;
wire      [7:0] XRAM_data_n1119;
wire      [7:0] XRAM_data_n1124;
wire      [7:0] XRAM_data_n1129;
wire      [7:0] XRAM_data_n1134;
wire      [7:0] XRAM_data_n1139;
wire      [7:0] XRAM_data_n1144;
wire      [7:0] XRAM_data_n1149;
wire      [7:0] XRAM_data_n1154;
wire      [7:0] XRAM_data_n1159;
wire      [7:0] XRAM_data_n1164;
wire      [7:0] XRAM_data_n1169;
wire      [7:0] XRAM_data_n1174;
wire      [7:0] XRAM_data_n1179;
wire      [7:0] XRAM_data_n1184;
wire      [7:0] XRAM_data_n1189;
wire      [7:0] XRAM_data_n1194;
wire      [7:0] XRAM_data_n1199;
wire      [7:0] XRAM_data_n1204;
wire      [7:0] XRAM_data_n1209;
wire      [7:0] XRAM_data_n1214;
wire      [7:0] XRAM_data_n1219;
wire      [7:0] XRAM_data_n1224;
wire      [7:0] XRAM_data_n1229;
wire      [7:0] XRAM_data_n915;
wire      [7:0] XRAM_data_n919;
wire      [7:0] XRAM_data_n924;
wire      [7:0] XRAM_data_n929;
wire      [7:0] XRAM_data_n934;
wire      [7:0] XRAM_data_n939;
wire      [7:0] XRAM_data_n944;
wire      [7:0] XRAM_data_n949;
wire      [7:0] XRAM_data_n954;
wire      [7:0] XRAM_data_n959;
wire      [7:0] XRAM_data_n964;
wire      [7:0] XRAM_data_n969;
wire      [7:0] XRAM_data_n974;
wire      [7:0] XRAM_data_n979;
wire      [7:0] XRAM_data_n984;
wire      [7:0] XRAM_data_n989;
wire      [7:0] XRAM_data_n994;
wire      [7:0] XRAM_data_n999;
wire            XRAM_wen0;
wire            XRAM_wen1;
wire            XRAM_wen2;
wire            XRAM_wen3;
wire            XRAM_wen4;
wire            XRAM_wen5;
wire            XRAM_wen6;
wire            XRAM_wen7;
wire    [159:0] __ILA_sha_acc_decode__;
wire            __ILA_sha_decode_of_I__DOT__0__;
wire            __ILA_sha_decode_of_I__DOT__100__;
wire            __ILA_sha_decode_of_I__DOT__101__;
wire            __ILA_sha_decode_of_I__DOT__102__;
wire            __ILA_sha_decode_of_I__DOT__103__;
wire            __ILA_sha_decode_of_I__DOT__104__;
wire            __ILA_sha_decode_of_I__DOT__105__;
wire            __ILA_sha_decode_of_I__DOT__106__;
wire            __ILA_sha_decode_of_I__DOT__107__;
wire            __ILA_sha_decode_of_I__DOT__108__;
wire            __ILA_sha_decode_of_I__DOT__109__;
wire            __ILA_sha_decode_of_I__DOT__10__;
wire            __ILA_sha_decode_of_I__DOT__110__;
wire            __ILA_sha_decode_of_I__DOT__111__;
wire            __ILA_sha_decode_of_I__DOT__112__;
wire            __ILA_sha_decode_of_I__DOT__113__;
wire            __ILA_sha_decode_of_I__DOT__114__;
wire            __ILA_sha_decode_of_I__DOT__115__;
wire            __ILA_sha_decode_of_I__DOT__116__;
wire            __ILA_sha_decode_of_I__DOT__117__;
wire            __ILA_sha_decode_of_I__DOT__118__;
wire            __ILA_sha_decode_of_I__DOT__119__;
wire            __ILA_sha_decode_of_I__DOT__11__;
wire            __ILA_sha_decode_of_I__DOT__120__;
wire            __ILA_sha_decode_of_I__DOT__121__;
wire            __ILA_sha_decode_of_I__DOT__122__;
wire            __ILA_sha_decode_of_I__DOT__123__;
wire            __ILA_sha_decode_of_I__DOT__124__;
wire            __ILA_sha_decode_of_I__DOT__125__;
wire            __ILA_sha_decode_of_I__DOT__126__;
wire            __ILA_sha_decode_of_I__DOT__127__;
wire            __ILA_sha_decode_of_I__DOT__128__;
wire            __ILA_sha_decode_of_I__DOT__129__;
wire            __ILA_sha_decode_of_I__DOT__12__;
wire            __ILA_sha_decode_of_I__DOT__130__;
wire            __ILA_sha_decode_of_I__DOT__131__;
wire            __ILA_sha_decode_of_I__DOT__132__;
wire            __ILA_sha_decode_of_I__DOT__133__;
wire            __ILA_sha_decode_of_I__DOT__134__;
wire            __ILA_sha_decode_of_I__DOT__135__;
wire            __ILA_sha_decode_of_I__DOT__136__;
wire            __ILA_sha_decode_of_I__DOT__137__;
wire            __ILA_sha_decode_of_I__DOT__138__;
wire            __ILA_sha_decode_of_I__DOT__139__;
wire            __ILA_sha_decode_of_I__DOT__13__;
wire            __ILA_sha_decode_of_I__DOT__140__;
wire            __ILA_sha_decode_of_I__DOT__141__;
wire            __ILA_sha_decode_of_I__DOT__142__;
wire            __ILA_sha_decode_of_I__DOT__143__;
wire            __ILA_sha_decode_of_I__DOT__144__;
wire            __ILA_sha_decode_of_I__DOT__145__;
wire            __ILA_sha_decode_of_I__DOT__146__;
wire            __ILA_sha_decode_of_I__DOT__147__;
wire            __ILA_sha_decode_of_I__DOT__148__;
wire            __ILA_sha_decode_of_I__DOT__149__;
wire            __ILA_sha_decode_of_I__DOT__14__;
wire            __ILA_sha_decode_of_I__DOT__150__;
wire            __ILA_sha_decode_of_I__DOT__151__;
wire            __ILA_sha_decode_of_I__DOT__152__;
wire            __ILA_sha_decode_of_I__DOT__153__;
wire            __ILA_sha_decode_of_I__DOT__154__;
wire            __ILA_sha_decode_of_I__DOT__155__;
wire            __ILA_sha_decode_of_I__DOT__156__;
wire            __ILA_sha_decode_of_I__DOT__157__;
wire            __ILA_sha_decode_of_I__DOT__158__;
wire            __ILA_sha_decode_of_I__DOT__159__;
wire            __ILA_sha_decode_of_I__DOT__15__;
wire            __ILA_sha_decode_of_I__DOT__16__;
wire            __ILA_sha_decode_of_I__DOT__17__;
wire            __ILA_sha_decode_of_I__DOT__18__;
wire            __ILA_sha_decode_of_I__DOT__19__;
wire            __ILA_sha_decode_of_I__DOT__1__;
wire            __ILA_sha_decode_of_I__DOT__20__;
wire            __ILA_sha_decode_of_I__DOT__21__;
wire            __ILA_sha_decode_of_I__DOT__22__;
wire            __ILA_sha_decode_of_I__DOT__23__;
wire            __ILA_sha_decode_of_I__DOT__24__;
wire            __ILA_sha_decode_of_I__DOT__25__;
wire            __ILA_sha_decode_of_I__DOT__26__;
wire            __ILA_sha_decode_of_I__DOT__27__;
wire            __ILA_sha_decode_of_I__DOT__28__;
wire            __ILA_sha_decode_of_I__DOT__29__;
wire            __ILA_sha_decode_of_I__DOT__2__;
wire            __ILA_sha_decode_of_I__DOT__30__;
wire            __ILA_sha_decode_of_I__DOT__31__;
wire            __ILA_sha_decode_of_I__DOT__32__;
wire            __ILA_sha_decode_of_I__DOT__33__;
wire            __ILA_sha_decode_of_I__DOT__34__;
wire            __ILA_sha_decode_of_I__DOT__35__;
wire            __ILA_sha_decode_of_I__DOT__36__;
wire            __ILA_sha_decode_of_I__DOT__37__;
wire            __ILA_sha_decode_of_I__DOT__38__;
wire            __ILA_sha_decode_of_I__DOT__39__;
wire            __ILA_sha_decode_of_I__DOT__3__;
wire            __ILA_sha_decode_of_I__DOT__40__;
wire            __ILA_sha_decode_of_I__DOT__41__;
wire            __ILA_sha_decode_of_I__DOT__42__;
wire            __ILA_sha_decode_of_I__DOT__43__;
wire            __ILA_sha_decode_of_I__DOT__44__;
wire            __ILA_sha_decode_of_I__DOT__45__;
wire            __ILA_sha_decode_of_I__DOT__46__;
wire            __ILA_sha_decode_of_I__DOT__47__;
wire            __ILA_sha_decode_of_I__DOT__48__;
wire            __ILA_sha_decode_of_I__DOT__49__;
wire            __ILA_sha_decode_of_I__DOT__4__;
wire            __ILA_sha_decode_of_I__DOT__50__;
wire            __ILA_sha_decode_of_I__DOT__51__;
wire            __ILA_sha_decode_of_I__DOT__52__;
wire            __ILA_sha_decode_of_I__DOT__53__;
wire            __ILA_sha_decode_of_I__DOT__54__;
wire            __ILA_sha_decode_of_I__DOT__55__;
wire            __ILA_sha_decode_of_I__DOT__56__;
wire            __ILA_sha_decode_of_I__DOT__57__;
wire            __ILA_sha_decode_of_I__DOT__58__;
wire            __ILA_sha_decode_of_I__DOT__59__;
wire            __ILA_sha_decode_of_I__DOT__5__;
wire            __ILA_sha_decode_of_I__DOT__60__;
wire            __ILA_sha_decode_of_I__DOT__61__;
wire            __ILA_sha_decode_of_I__DOT__62__;
wire            __ILA_sha_decode_of_I__DOT__63__;
wire            __ILA_sha_decode_of_I__DOT__64__;
wire            __ILA_sha_decode_of_I__DOT__65__;
wire            __ILA_sha_decode_of_I__DOT__66__;
wire            __ILA_sha_decode_of_I__DOT__67__;
wire            __ILA_sha_decode_of_I__DOT__68__;
wire            __ILA_sha_decode_of_I__DOT__69__;
wire            __ILA_sha_decode_of_I__DOT__6__;
wire            __ILA_sha_decode_of_I__DOT__70__;
wire            __ILA_sha_decode_of_I__DOT__71__;
wire            __ILA_sha_decode_of_I__DOT__72__;
wire            __ILA_sha_decode_of_I__DOT__73__;
wire            __ILA_sha_decode_of_I__DOT__74__;
wire            __ILA_sha_decode_of_I__DOT__75__;
wire            __ILA_sha_decode_of_I__DOT__76__;
wire            __ILA_sha_decode_of_I__DOT__77__;
wire            __ILA_sha_decode_of_I__DOT__78__;
wire            __ILA_sha_decode_of_I__DOT__79__;
wire            __ILA_sha_decode_of_I__DOT__7__;
wire            __ILA_sha_decode_of_I__DOT__80__;
wire            __ILA_sha_decode_of_I__DOT__81__;
wire            __ILA_sha_decode_of_I__DOT__82__;
wire            __ILA_sha_decode_of_I__DOT__83__;
wire            __ILA_sha_decode_of_I__DOT__84__;
wire            __ILA_sha_decode_of_I__DOT__85__;
wire            __ILA_sha_decode_of_I__DOT__86__;
wire            __ILA_sha_decode_of_I__DOT__87__;
wire            __ILA_sha_decode_of_I__DOT__88__;
wire            __ILA_sha_decode_of_I__DOT__89__;
wire            __ILA_sha_decode_of_I__DOT__8__;
wire            __ILA_sha_decode_of_I__DOT__90__;
wire            __ILA_sha_decode_of_I__DOT__91__;
wire            __ILA_sha_decode_of_I__DOT__92__;
wire            __ILA_sha_decode_of_I__DOT__93__;
wire            __ILA_sha_decode_of_I__DOT__94__;
wire            __ILA_sha_decode_of_I__DOT__95__;
wire            __ILA_sha_decode_of_I__DOT__96__;
wire            __ILA_sha_decode_of_I__DOT__97__;
wire            __ILA_sha_decode_of_I__DOT__98__;
wire            __ILA_sha_decode_of_I__DOT__99__;
wire            __ILA_sha_decode_of_I__DOT__9__;
wire    [159:0] __ILA_sha_grant__;
wire            __ILA_sha_valid__;
wire            clk;
wire      [1:0] cmd;
wire     [15:0] cmdaddr;
wire      [7:0] cmddata;
wire            n0;
wire            n1;
wire            n10;
wire            n100;
wire      [7:0] n1000;
wire    [143:0] n1001;
wire     [15:0] n1002;
wire      [7:0] n1005;
wire    [151:0] n1006;
wire     [15:0] n1007;
wire            n101;
wire      [7:0] n1010;
wire    [159:0] n1011;
wire     [15:0] n1012;
wire      [7:0] n1015;
wire    [167:0] n1016;
wire     [15:0] n1017;
wire            n102;
wire      [7:0] n1020;
wire    [175:0] n1021;
wire     [15:0] n1022;
wire      [7:0] n1025;
wire    [183:0] n1026;
wire     [15:0] n1027;
wire            n103;
wire      [7:0] n1030;
wire    [191:0] n1031;
wire     [15:0] n1032;
wire      [7:0] n1035;
wire    [199:0] n1036;
wire     [15:0] n1037;
wire            n104;
wire      [7:0] n1040;
wire    [207:0] n1041;
wire     [15:0] n1042;
wire      [7:0] n1045;
wire    [215:0] n1046;
wire     [15:0] n1047;
wire            n105;
wire      [7:0] n1050;
wire    [223:0] n1051;
wire     [15:0] n1052;
wire      [7:0] n1055;
wire    [231:0] n1056;
wire     [15:0] n1057;
wire            n106;
wire      [7:0] n1060;
wire    [239:0] n1061;
wire     [15:0] n1062;
wire      [7:0] n1065;
wire    [247:0] n1066;
wire     [15:0] n1067;
wire            n107;
wire      [7:0] n1070;
wire    [255:0] n1071;
wire     [15:0] n1072;
wire      [7:0] n1075;
wire    [263:0] n1076;
wire     [15:0] n1077;
wire            n108;
wire      [7:0] n1080;
wire    [271:0] n1081;
wire     [15:0] n1082;
wire      [7:0] n1085;
wire    [279:0] n1086;
wire     [15:0] n1087;
wire            n109;
wire      [7:0] n1090;
wire    [287:0] n1091;
wire     [15:0] n1092;
wire      [7:0] n1095;
wire    [295:0] n1096;
wire     [15:0] n1097;
wire            n11;
wire            n110;
wire      [7:0] n1100;
wire    [303:0] n1101;
wire     [15:0] n1102;
wire      [7:0] n1105;
wire    [311:0] n1106;
wire     [15:0] n1107;
wire            n111;
wire      [7:0] n1110;
wire    [319:0] n1111;
wire     [15:0] n1112;
wire      [7:0] n1115;
wire    [327:0] n1116;
wire     [15:0] n1117;
wire            n112;
wire      [7:0] n1120;
wire    [335:0] n1121;
wire     [15:0] n1122;
wire      [7:0] n1125;
wire    [343:0] n1126;
wire     [15:0] n1127;
wire            n113;
wire      [7:0] n1130;
wire    [351:0] n1131;
wire     [15:0] n1132;
wire      [7:0] n1135;
wire    [359:0] n1136;
wire     [15:0] n1137;
wire            n114;
wire      [7:0] n1140;
wire    [367:0] n1141;
wire     [15:0] n1142;
wire      [7:0] n1145;
wire    [375:0] n1146;
wire     [15:0] n1147;
wire            n115;
wire      [7:0] n1150;
wire    [383:0] n1151;
wire     [15:0] n1152;
wire      [7:0] n1155;
wire    [391:0] n1156;
wire     [15:0] n1157;
wire            n116;
wire      [7:0] n1160;
wire    [399:0] n1161;
wire     [15:0] n1162;
wire      [7:0] n1165;
wire    [407:0] n1166;
wire     [15:0] n1167;
wire            n117;
wire      [7:0] n1170;
wire    [415:0] n1171;
wire     [15:0] n1172;
wire      [7:0] n1175;
wire    [423:0] n1176;
wire     [15:0] n1177;
wire            n118;
wire      [7:0] n1180;
wire    [431:0] n1181;
wire     [15:0] n1182;
wire      [7:0] n1185;
wire    [439:0] n1186;
wire     [15:0] n1187;
wire            n119;
wire      [7:0] n1190;
wire    [447:0] n1191;
wire     [15:0] n1192;
wire      [7:0] n1195;
wire    [455:0] n1196;
wire     [15:0] n1197;
wire            n12;
wire            n120;
wire      [7:0] n1200;
wire    [463:0] n1201;
wire     [15:0] n1202;
wire      [7:0] n1205;
wire    [471:0] n1206;
wire     [15:0] n1207;
wire            n121;
wire      [7:0] n1210;
wire    [479:0] n1211;
wire     [15:0] n1212;
wire      [7:0] n1215;
wire    [487:0] n1216;
wire     [15:0] n1217;
wire            n122;
wire      [7:0] n1220;
wire    [495:0] n1221;
wire     [15:0] n1222;
wire      [7:0] n1225;
wire    [503:0] n1226;
wire     [15:0] n1227;
wire            n123;
wire      [7:0] n1230;
wire    [511:0] n1231;
wire    [511:0] n1232;
wire      [7:0] n1233;
wire     [15:0] n1234;
wire      [7:0] n1235;
wire     [15:0] n1236;
wire            n1237;
wire            n1238;
wire            n1239;
wire            n124;
wire            n1240;
wire            n1241;
wire            n1242;
wire            n1243;
wire            n1244;
wire            n1245;
wire            n1246;
wire            n1247;
wire            n1248;
wire            n1249;
wire            n125;
wire            n1250;
wire            n1251;
wire            n1252;
wire            n1253;
wire            n1254;
wire            n1255;
wire            n1256;
wire            n1257;
wire            n1258;
wire            n1259;
wire            n126;
wire            n1260;
wire            n1261;
wire            n1262;
wire            n1263;
wire            n1264;
wire            n1265;
wire            n1266;
wire            n1267;
wire            n1268;
wire            n1269;
wire            n127;
wire            n1270;
wire            n1271;
wire            n1272;
wire            n1273;
wire            n1274;
wire            n1275;
wire            n1276;
wire            n1277;
wire            n1278;
wire            n1279;
wire            n128;
wire            n1280;
wire            n1281;
wire            n1282;
wire            n1283;
wire            n1284;
wire            n1285;
wire            n1286;
wire            n1287;
wire            n1288;
wire            n1289;
wire            n129;
wire            n1290;
wire            n1291;
wire            n1292;
wire            n1293;
wire            n1294;
wire            n1295;
wire            n1296;
wire            n1297;
wire            n1298;
wire            n1299;
wire            n13;
wire            n130;
wire            n1300;
wire            n1301;
wire            n1302;
wire            n1303;
wire            n1304;
wire            n1305;
wire            n1306;
wire            n1307;
wire            n1308;
wire            n1309;
wire            n131;
wire            n1310;
wire            n1311;
wire            n1312;
wire            n1313;
wire            n1314;
wire            n1315;
wire            n1316;
wire            n1317;
wire            n1318;
wire      [2:0] n1319;
wire            n132;
wire            n1320;
wire            n1321;
wire            n1322;
wire            n1323;
wire            n1324;
wire            n1325;
wire            n1326;
wire            n1327;
wire            n1328;
wire            n1329;
wire            n133;
wire            n1330;
wire            n1331;
wire            n1332;
wire            n1333;
wire            n1334;
wire            n1335;
wire            n1336;
wire            n1337;
wire            n1338;
wire            n1339;
wire            n134;
wire            n1340;
wire            n1341;
wire            n1342;
wire            n1343;
wire            n1344;
wire            n1345;
wire            n1346;
wire            n1347;
wire            n1348;
wire            n1349;
wire            n135;
wire            n1350;
wire            n1351;
wire            n1352;
wire            n1353;
wire            n1354;
wire            n1355;
wire            n1356;
wire            n1357;
wire            n1358;
wire            n1359;
wire            n136;
wire            n1360;
wire            n1361;
wire            n1362;
wire            n1363;
wire            n1364;
wire            n1365;
wire            n1366;
wire            n1367;
wire            n1368;
wire            n1369;
wire            n137;
wire            n1370;
wire            n1371;
wire            n1372;
wire            n1373;
wire            n1374;
wire            n1375;
wire            n1376;
wire            n1377;
wire            n1378;
wire            n1379;
wire            n138;
wire            n1380;
wire            n1381;
wire            n1382;
wire            n1383;
wire            n1384;
wire            n1385;
wire            n1386;
wire            n1387;
wire            n1388;
wire            n1389;
wire            n139;
wire            n1390;
wire            n1391;
wire            n1392;
wire            n1393;
wire            n1394;
wire            n1395;
wire            n1396;
wire            n1397;
wire            n1398;
wire            n1399;
wire            n14;
wire            n140;
wire            n1400;
wire            n1401;
wire            n1402;
wire            n1403;
wire            n1404;
wire            n1405;
wire            n1406;
wire            n1407;
wire            n1408;
wire            n1409;
wire            n141;
wire            n1410;
wire            n1411;
wire            n1412;
wire            n1413;
wire            n1414;
wire            n1415;
wire            n1416;
wire            n1417;
wire            n1418;
wire            n1419;
wire            n142;
wire            n1420;
wire            n1421;
wire            n1422;
wire            n1423;
wire            n1424;
wire            n1425;
wire            n1426;
wire            n1427;
wire            n1428;
wire            n1429;
wire            n143;
wire            n1430;
wire            n1431;
wire            n1432;
wire            n1433;
wire            n1434;
wire            n1435;
wire            n1436;
wire            n1437;
wire            n1438;
wire            n1439;
wire            n144;
wire            n1440;
wire            n1441;
wire            n1442;
wire            n1443;
wire            n1444;
wire            n1445;
wire            n1446;
wire            n1447;
wire            n1448;
wire            n1449;
wire            n145;
wire            n1450;
wire            n1451;
wire            n1452;
wire            n1453;
wire            n1454;
wire            n1455;
wire            n1456;
wire            n1457;
wire            n1458;
wire            n1459;
wire            n146;
wire            n1460;
wire            n1461;
wire            n1462;
wire            n1463;
wire            n1464;
wire            n1465;
wire            n1466;
wire            n1467;
wire            n1468;
wire            n1469;
wire            n147;
wire            n1470;
wire            n1471;
wire            n1472;
wire            n1473;
wire            n1474;
wire            n1475;
wire            n1476;
wire            n1477;
wire            n1478;
wire            n1479;
wire            n148;
wire            n1480;
wire            n1481;
wire            n1482;
wire            n1483;
wire            n1484;
wire            n1485;
wire            n1486;
wire            n1487;
wire            n1488;
wire            n1489;
wire            n149;
wire            n1490;
wire            n1491;
wire            n1492;
wire            n1493;
wire            n1494;
wire            n1495;
wire            n1496;
wire            n1497;
wire            n1498;
wire            n1499;
wire            n15;
wire            n150;
wire            n1500;
wire            n1501;
wire            n1502;
wire            n1503;
wire            n1504;
wire            n1505;
wire            n1506;
wire            n1507;
wire            n1508;
wire            n1509;
wire            n151;
wire            n1510;
wire            n1511;
wire            n1512;
wire            n1513;
wire            n1514;
wire            n1515;
wire            n1516;
wire            n1517;
wire            n1518;
wire            n1519;
wire            n152;
wire            n1520;
wire            n1521;
wire            n1522;
wire            n1523;
wire            n1524;
wire            n1525;
wire            n1526;
wire            n1527;
wire            n1528;
wire            n1529;
wire            n153;
wire            n1530;
wire            n1531;
wire            n1532;
wire            n1533;
wire            n1534;
wire            n1535;
wire            n1536;
wire            n1537;
wire            n1538;
wire            n1539;
wire            n154;
wire            n1540;
wire            n1541;
wire            n1542;
wire            n1543;
wire            n1544;
wire            n1545;
wire            n1546;
wire            n1547;
wire            n1548;
wire            n1549;
wire            n155;
wire            n1550;
wire            n1551;
wire            n1552;
wire            n1553;
wire            n1554;
wire            n1555;
wire            n1556;
wire            n1557;
wire            n1558;
wire            n1559;
wire            n156;
wire            n1560;
wire            n1561;
wire            n1562;
wire            n1563;
wire            n1564;
wire            n1565;
wire            n1566;
wire            n1567;
wire            n1568;
wire            n1569;
wire            n157;
wire            n1570;
wire            n1571;
wire            n1572;
wire            n1573;
wire            n1574;
wire            n1575;
wire            n1576;
wire            n1577;
wire            n1578;
wire            n1579;
wire            n158;
wire            n1580;
wire            n1581;
wire            n1582;
wire            n1583;
wire            n1584;
wire            n1585;
wire            n1586;
wire            n1587;
wire            n1588;
wire            n1589;
wire            n159;
wire            n1590;
wire            n1591;
wire            n1592;
wire            n1593;
wire            n1594;
wire            n1595;
wire            n1596;
wire            n1597;
wire            n1598;
wire            n1599;
wire            n16;
wire            n160;
wire            n1600;
wire            n1601;
wire            n1602;
wire            n1603;
wire            n1604;
wire            n1605;
wire            n1606;
wire            n1607;
wire            n1608;
wire            n1609;
wire            n161;
wire            n1610;
wire            n1611;
wire            n1612;
wire            n1613;
wire            n1614;
wire            n1615;
wire            n1616;
wire            n1617;
wire            n1618;
wire            n1619;
wire            n162;
wire            n1620;
wire            n1621;
wire            n1622;
wire            n1623;
wire            n1624;
wire            n1625;
wire            n1626;
wire            n1627;
wire            n1628;
wire      [2:0] n1629;
wire            n163;
wire      [2:0] n1630;
wire      [2:0] n1631;
wire      [2:0] n1632;
wire            n1633;
wire      [2:0] n1634;
wire      [7:0] n1635;
wire     [15:0] n1636;
wire      [7:0] n1637;
wire     [15:0] n1638;
wire            n1639;
wire            n164;
wire            n1640;
wire            n1641;
wire            n1642;
wire            n1643;
wire            n1644;
wire            n1645;
wire            n1646;
wire            n1647;
wire            n1648;
wire            n1649;
wire            n165;
wire            n1650;
wire            n1651;
wire            n1652;
wire            n1653;
wire            n1654;
wire            n1655;
wire            n1656;
wire            n1657;
wire            n1658;
wire            n1659;
wire            n166;
wire            n1660;
wire            n1661;
wire            n1662;
wire            n1663;
wire            n1664;
wire            n1665;
wire            n1666;
wire            n1667;
wire            n1668;
wire            n1669;
wire            n167;
wire            n1670;
wire            n1671;
wire            n1672;
wire            n1673;
wire            n1674;
wire            n1675;
wire            n1676;
wire            n1677;
wire            n1678;
wire            n1679;
wire            n168;
wire            n1680;
wire            n1681;
wire            n1682;
wire            n1683;
wire            n1684;
wire            n1685;
wire            n1686;
wire            n1687;
wire            n1688;
wire            n1689;
wire            n169;
wire            n1690;
wire            n1691;
wire            n1692;
wire            n1693;
wire            n1694;
wire            n1695;
wire            n1696;
wire            n1697;
wire            n1698;
wire            n1699;
wire            n17;
wire            n170;
wire            n1700;
wire            n1701;
wire            n1702;
wire            n1703;
wire            n1704;
wire            n1705;
wire            n1706;
wire            n1707;
wire            n1708;
wire            n1709;
wire            n171;
wire            n1710;
wire            n1711;
wire            n1712;
wire            n1713;
wire            n1714;
wire            n1715;
wire            n1716;
wire            n1717;
wire            n1718;
wire            n1719;
wire            n172;
wire            n1720;
wire            n1721;
wire            n1722;
wire            n1723;
wire            n1724;
wire            n1725;
wire            n1726;
wire            n1727;
wire            n1728;
wire            n1729;
wire            n173;
wire            n1730;
wire            n1731;
wire            n1732;
wire            n1733;
wire            n1734;
wire            n1735;
wire            n1736;
wire            n1737;
wire            n1738;
wire            n1739;
wire            n174;
wire            n1740;
wire            n1741;
wire            n1742;
wire            n1743;
wire            n1744;
wire            n1745;
wire            n1746;
wire            n1747;
wire            n1748;
wire            n1749;
wire            n175;
wire            n1750;
wire            n1751;
wire            n1752;
wire            n1753;
wire            n1754;
wire            n1755;
wire            n1756;
wire            n1757;
wire            n1758;
wire            n1759;
wire            n176;
wire            n1760;
wire            n1761;
wire            n1762;
wire            n1763;
wire            n1764;
wire            n1765;
wire            n1766;
wire            n1767;
wire            n1768;
wire            n1769;
wire            n177;
wire            n1770;
wire            n1771;
wire            n1772;
wire            n1773;
wire            n1774;
wire            n1775;
wire            n1776;
wire            n1777;
wire            n1778;
wire            n1779;
wire            n178;
wire            n1780;
wire            n1781;
wire            n1782;
wire            n1783;
wire            n1784;
wire            n1785;
wire            n1786;
wire            n1787;
wire            n1788;
wire            n1789;
wire            n179;
wire            n1790;
wire            n1791;
wire            n1792;
wire            n1793;
wire            n1794;
wire            n1795;
wire            n1796;
wire            n1797;
wire            n1798;
wire            n1799;
wire            n18;
wire            n180;
wire            n1800;
wire            n1801;
wire            n1802;
wire            n1803;
wire            n1804;
wire            n1805;
wire            n1806;
wire            n1807;
wire            n1808;
wire            n1809;
wire            n181;
wire            n1810;
wire            n1811;
wire            n1812;
wire            n1813;
wire            n1814;
wire            n1815;
wire            n1816;
wire            n1817;
wire            n1818;
wire            n1819;
wire            n182;
wire            n1820;
wire            n1821;
wire            n1822;
wire            n1823;
wire            n1824;
wire            n1825;
wire            n1826;
wire            n1827;
wire            n1828;
wire            n1829;
wire            n183;
wire            n1830;
wire            n1831;
wire            n1832;
wire            n1833;
wire            n1834;
wire            n1835;
wire            n1836;
wire            n1837;
wire            n1838;
wire            n1839;
wire            n184;
wire            n1840;
wire            n1841;
wire            n1842;
wire            n1843;
wire            n1844;
wire            n1845;
wire            n1846;
wire            n1847;
wire            n1848;
wire            n1849;
wire            n185;
wire            n1850;
wire            n1851;
wire            n1852;
wire            n1853;
wire            n1854;
wire            n1855;
wire            n1856;
wire            n1857;
wire            n1858;
wire            n1859;
wire            n186;
wire            n1860;
wire            n1861;
wire            n1862;
wire            n1863;
wire            n1864;
wire            n1865;
wire            n1866;
wire            n1867;
wire            n1868;
wire            n1869;
wire            n187;
wire            n1870;
wire            n1871;
wire            n1872;
wire            n1873;
wire            n1874;
wire            n1875;
wire            n1876;
wire            n1877;
wire            n1878;
wire            n1879;
wire            n188;
wire            n1880;
wire            n1881;
wire            n1882;
wire            n1883;
wire            n1884;
wire            n1885;
wire            n1886;
wire            n1887;
wire            n1888;
wire            n1889;
wire            n189;
wire            n1890;
wire            n1891;
wire            n1892;
wire            n1893;
wire            n1894;
wire            n1895;
wire            n1896;
wire            n1897;
wire            n1898;
wire            n1899;
wire            n19;
wire            n190;
wire            n1900;
wire            n1901;
wire            n1902;
wire            n1903;
wire            n1904;
wire            n1905;
wire            n1906;
wire            n1907;
wire            n1908;
wire            n1909;
wire            n191;
wire            n1910;
wire            n1911;
wire            n1912;
wire            n1913;
wire            n1914;
wire            n1915;
wire            n1916;
wire            n1917;
wire            n1918;
wire            n1919;
wire            n192;
wire            n1920;
wire            n1921;
wire            n1922;
wire            n1923;
wire            n1924;
wire            n1925;
wire            n1926;
wire            n1927;
wire            n1928;
wire            n1929;
wire            n193;
wire            n1930;
wire            n1931;
wire            n1932;
wire            n1933;
wire            n1934;
wire            n1935;
wire            n1936;
wire            n1937;
wire            n1938;
wire            n1939;
wire            n194;
wire            n1940;
wire            n1941;
wire            n1942;
wire            n1943;
wire            n1944;
wire            n1945;
wire            n1946;
wire            n1947;
wire            n1948;
wire            n1949;
wire            n195;
wire            n1950;
wire            n1951;
wire            n1952;
wire            n1953;
wire            n1954;
wire            n1955;
wire            n1956;
wire            n1957;
wire            n1958;
wire            n1959;
wire            n196;
wire            n1960;
wire            n1961;
wire            n1962;
wire            n1963;
wire            n1964;
wire            n1965;
wire            n1966;
wire            n1967;
wire            n1968;
wire            n1969;
wire            n197;
wire            n1970;
wire            n1971;
wire            n1972;
wire            n1973;
wire            n1974;
wire            n1975;
wire            n1976;
wire            n1977;
wire            n1978;
wire            n1979;
wire            n198;
wire            n1980;
wire            n1981;
wire            n1982;
wire            n1983;
wire            n1984;
wire            n1985;
wire            n1986;
wire            n1987;
wire            n1988;
wire            n1989;
wire            n199;
wire            n1990;
wire            n1991;
wire            n1992;
wire            n1993;
wire            n1994;
wire            n1995;
wire            n1996;
wire            n1997;
wire            n1998;
wire            n1999;
wire            n2;
wire            n20;
wire            n200;
wire            n2000;
wire            n2001;
wire            n2002;
wire            n2003;
wire            n2004;
wire            n2005;
wire            n2006;
wire            n2007;
wire            n2008;
wire            n2009;
wire            n201;
wire            n2010;
wire            n2011;
wire            n2012;
wire            n2013;
wire            n2014;
wire            n2015;
wire            n2016;
wire            n2017;
wire            n2018;
wire            n2019;
wire            n202;
wire            n2020;
wire            n2021;
wire            n2022;
wire            n2023;
wire            n2024;
wire            n2025;
wire            n2026;
wire            n2027;
wire            n2028;
wire            n2029;
wire            n203;
wire            n2030;
wire            n2031;
wire            n2032;
wire            n2033;
wire            n2034;
wire            n2035;
wire            n2036;
wire            n2037;
wire            n2038;
wire            n2039;
wire            n204;
wire            n2040;
wire            n2041;
wire            n2042;
wire            n2043;
wire            n2044;
wire            n2045;
wire            n2046;
wire            n2047;
wire            n2048;
wire            n2049;
wire            n205;
wire            n2050;
wire            n2051;
wire            n2052;
wire            n2053;
wire            n2054;
wire            n2055;
wire            n2056;
wire            n2057;
wire            n2058;
wire            n2059;
wire            n206;
wire            n2060;
wire            n2061;
wire            n2062;
wire            n2063;
wire            n2064;
wire            n2065;
wire            n2066;
wire            n2067;
wire            n2068;
wire            n2069;
wire            n207;
wire            n2070;
wire            n2071;
wire            n2072;
wire            n2073;
wire            n2074;
wire            n2075;
wire            n2076;
wire            n2077;
wire            n2078;
wire            n2079;
wire            n208;
wire            n2080;
wire            n2081;
wire            n2082;
wire            n2083;
wire            n2084;
wire            n2085;
wire            n2086;
wire            n2087;
wire            n2088;
wire            n2089;
wire            n209;
wire            n2090;
wire            n2091;
wire            n2092;
wire            n2093;
wire            n2094;
wire            n2095;
wire            n2096;
wire            n2097;
wire            n2098;
wire            n2099;
wire            n21;
wire            n210;
wire            n2100;
wire            n2101;
wire            n2102;
wire            n2103;
wire            n2104;
wire            n2105;
wire            n2106;
wire            n2107;
wire            n2108;
wire            n2109;
wire            n211;
wire            n2110;
wire            n2111;
wire            n2112;
wire            n2113;
wire            n2114;
wire            n2115;
wire            n2116;
wire            n2117;
wire            n2118;
wire            n2119;
wire            n212;
wire            n2120;
wire            n2121;
wire            n2122;
wire            n2123;
wire            n2124;
wire            n2125;
wire            n2126;
wire            n2127;
wire            n2128;
wire            n2129;
wire            n213;
wire            n2130;
wire            n2131;
wire            n2132;
wire            n2133;
wire            n2134;
wire            n2135;
wire            n2136;
wire            n2137;
wire            n2138;
wire            n2139;
wire            n214;
wire            n2140;
wire            n2141;
wire            n2142;
wire            n2143;
wire            n2144;
wire            n2145;
wire            n2146;
wire            n2147;
wire            n2148;
wire            n2149;
wire            n215;
wire            n2150;
wire            n2151;
wire            n2152;
wire            n2153;
wire            n2154;
wire            n2155;
wire            n2156;
wire            n2157;
wire            n2158;
wire            n2159;
wire            n216;
wire            n2160;
wire            n2161;
wire            n2162;
wire            n2163;
wire            n2164;
wire            n2165;
wire            n2166;
wire            n2167;
wire            n2168;
wire            n2169;
wire            n217;
wire            n2170;
wire            n2171;
wire            n2172;
wire            n2173;
wire            n2174;
wire            n2175;
wire            n2176;
wire            n2177;
wire            n2178;
wire            n2179;
wire      [7:0] n218;
wire            n2180;
wire            n2181;
wire            n2182;
wire            n2183;
wire            n2184;
wire            n2185;
wire            n2186;
wire            n2187;
wire            n2188;
wire            n2189;
wire            n219;
wire            n2190;
wire            n2191;
wire            n2192;
wire            n2193;
wire            n2194;
wire            n2195;
wire            n2196;
wire            n2197;
wire            n2198;
wire            n2199;
wire            n22;
wire            n220;
wire            n2200;
wire            n2201;
wire            n2202;
wire            n2203;
wire            n2204;
wire            n2205;
wire            n2206;
wire            n2207;
wire            n2208;
wire            n2209;
wire            n221;
wire            n2210;
wire            n2211;
wire            n2212;
wire            n2213;
wire            n2214;
wire            n2215;
wire            n2216;
wire            n2217;
wire            n2218;
wire            n2219;
wire            n222;
wire            n2220;
wire            n2221;
wire            n2222;
wire            n2223;
wire            n2224;
wire            n2225;
wire            n2226;
wire            n2227;
wire            n2228;
wire            n2229;
wire            n223;
wire            n2230;
wire            n2231;
wire            n2232;
wire            n2233;
wire            n2234;
wire            n2235;
wire            n2236;
wire            n2237;
wire            n2238;
wire            n2239;
wire            n224;
wire            n2240;
wire            n2241;
wire            n2242;
wire            n2243;
wire            n2244;
wire            n2245;
wire            n2246;
wire            n2247;
wire            n2248;
wire            n2249;
wire            n225;
wire            n2250;
wire            n2251;
wire            n2252;
wire            n2253;
wire            n2254;
wire            n2255;
wire            n2256;
wire            n2257;
wire            n2258;
wire            n2259;
wire            n226;
wire            n2260;
wire            n2261;
wire            n2262;
wire            n2263;
wire            n2264;
wire            n2265;
wire            n2266;
wire            n2267;
wire            n2268;
wire            n2269;
wire            n227;
wire            n2270;
wire            n2271;
wire            n2272;
wire            n2273;
wire            n2274;
wire            n2275;
wire            n2276;
wire            n2277;
wire            n2278;
wire            n2279;
wire            n228;
wire            n2280;
wire            n2281;
wire            n2282;
wire            n2283;
wire            n2284;
wire            n2285;
wire            n2286;
wire            n2287;
wire            n2288;
wire            n2289;
wire            n229;
wire            n2290;
wire            n2291;
wire            n2292;
wire            n2293;
wire            n2294;
wire            n2295;
wire            n2296;
wire            n2297;
wire            n2298;
wire            n2299;
wire            n23;
wire            n230;
wire            n2300;
wire            n2301;
wire            n2302;
wire            n2303;
wire            n2304;
wire            n2305;
wire            n2306;
wire            n2307;
wire            n2308;
wire            n2309;
wire            n231;
wire            n2310;
wire            n2311;
wire            n2312;
wire            n2313;
wire            n2314;
wire            n2315;
wire            n2316;
wire            n2317;
wire            n2318;
wire            n2319;
wire            n232;
wire            n2320;
wire            n2321;
wire            n2322;
wire            n2323;
wire            n2324;
wire            n2325;
wire            n2326;
wire            n2327;
wire            n2328;
wire            n2329;
wire            n233;
wire            n2330;
wire            n2331;
wire            n2332;
wire            n2333;
wire            n2334;
wire            n2335;
wire            n2336;
wire            n2337;
wire            n2338;
wire            n2339;
wire            n234;
wire            n2340;
wire            n2341;
wire            n2342;
wire            n2343;
wire            n2344;
wire            n2345;
wire            n2346;
wire            n2347;
wire            n2348;
wire            n2349;
wire            n235;
wire            n2350;
wire            n2351;
wire            n2352;
wire            n2353;
wire            n2354;
wire            n2355;
wire            n2356;
wire            n2357;
wire            n2358;
wire            n2359;
wire            n236;
wire            n2360;
wire            n2361;
wire            n2362;
wire            n2363;
wire            n2364;
wire            n2365;
wire     [15:0] n2366;
wire      [7:0] n2367;
wire     [15:0] n2368;
wire      [7:0] n2369;
wire            n237;
wire     [15:0] n2370;
wire      [7:0] n2371;
wire     [15:0] n2372;
wire      [7:0] n2373;
wire     [15:0] n2374;
wire      [7:0] n2375;
wire     [15:0] n2376;
wire      [7:0] n2377;
wire     [15:0] n2378;
wire      [7:0] n2379;
wire            n238;
wire     [15:0] n2380;
wire      [7:0] n2381;
wire            n2382;
wire            n2383;
wire            n2384;
wire            n2385;
wire            n2386;
wire            n2387;
wire            n2388;
wire            n2389;
wire            n239;
wire            n2390;
wire            n2391;
wire            n2392;
wire            n2393;
wire            n2394;
wire            n2395;
wire            n2396;
wire            n2397;
wire            n2398;
wire            n2399;
wire            n24;
wire      [7:0] n240;
wire            n2400;
wire            n2401;
wire            n2402;
wire            n2403;
wire            n2404;
wire            n2405;
wire            n2406;
wire            n2407;
wire            n2408;
wire            n2409;
wire            n241;
wire            n2410;
wire            n2411;
wire            n2412;
wire            n2413;
wire            n2414;
wire            n2415;
wire            n2416;
wire            n2417;
wire            n2418;
wire            n2419;
wire            n242;
wire            n2420;
wire            n2421;
wire            n2422;
wire            n2423;
wire            n2424;
wire            n2425;
wire            n2426;
wire            n2427;
wire            n2428;
wire            n2429;
wire            n243;
wire            n2430;
wire            n2431;
wire            n2432;
wire            n2433;
wire            n2434;
wire            n2435;
wire            n2436;
wire            n2437;
wire            n2438;
wire            n2439;
wire            n244;
wire            n2440;
wire            n2441;
wire            n2442;
wire            n2443;
wire            n2444;
wire            n2445;
wire            n2446;
wire            n2447;
wire            n2448;
wire            n2449;
wire            n245;
wire            n2450;
wire            n2451;
wire            n2452;
wire            n2453;
wire            n2454;
wire            n2455;
wire            n2456;
wire            n2457;
wire            n2458;
wire            n2459;
wire            n246;
wire            n2460;
wire            n2461;
wire            n2462;
wire            n2463;
wire            n2464;
wire            n2465;
wire            n2466;
wire            n2467;
wire            n2468;
wire            n2469;
wire            n247;
wire            n2470;
wire            n2471;
wire            n2472;
wire            n2473;
wire            n2474;
wire            n2475;
wire            n2476;
wire            n2477;
wire            n2478;
wire            n2479;
wire            n248;
wire            n2480;
wire            n2481;
wire            n2482;
wire            n2483;
wire            n2484;
wire            n2485;
wire            n2486;
wire            n2487;
wire            n2488;
wire            n2489;
wire            n249;
wire            n2490;
wire            n2491;
wire            n2492;
wire            n2493;
wire            n2494;
wire            n2495;
wire            n2496;
wire            n2497;
wire            n2498;
wire            n2499;
wire            n25;
wire            n250;
wire            n2500;
wire            n2501;
wire            n2502;
wire            n2503;
wire            n2504;
wire            n2505;
wire            n2506;
wire            n2507;
wire            n2508;
wire            n2509;
wire            n251;
wire            n2510;
wire            n2511;
wire            n2512;
wire            n2513;
wire            n2514;
wire            n2515;
wire            n2516;
wire            n2517;
wire            n2518;
wire            n2519;
wire            n252;
wire            n2520;
wire            n2521;
wire            n2522;
wire            n2523;
wire            n2524;
wire            n2525;
wire            n2526;
wire            n2527;
wire            n2528;
wire            n2529;
wire            n253;
wire            n2530;
wire            n2531;
wire            n2532;
wire            n2533;
wire            n2534;
wire            n2535;
wire            n2536;
wire            n2537;
wire            n2538;
wire            n2539;
wire            n254;
wire            n2540;
wire            n2541;
wire            n2542;
wire            n2543;
wire            n2544;
wire            n2545;
wire            n2546;
wire            n2547;
wire            n2548;
wire            n2549;
wire            n255;
wire            n2550;
wire            n2551;
wire            n2552;
wire            n2553;
wire            n2554;
wire            n2555;
wire            n2556;
wire            n2557;
wire            n2558;
wire            n2559;
wire            n256;
wire            n2560;
wire            n2561;
wire            n2562;
wire            n2563;
wire            n2564;
wire            n2565;
wire            n2566;
wire            n2567;
wire            n2568;
wire            n2569;
wire            n257;
wire            n2570;
wire            n2571;
wire            n2572;
wire            n2573;
wire            n2574;
wire            n2575;
wire            n2576;
wire            n2577;
wire            n2578;
wire            n2579;
wire            n258;
wire            n2580;
wire            n2581;
wire            n2582;
wire            n2583;
wire            n2584;
wire            n2585;
wire            n2586;
wire            n2587;
wire            n2588;
wire            n2589;
wire            n259;
wire            n2590;
wire            n2591;
wire            n2592;
wire            n2593;
wire            n2594;
wire            n2595;
wire            n2596;
wire            n2597;
wire            n2598;
wire            n2599;
wire            n26;
wire            n260;
wire            n2600;
wire            n2601;
wire            n2602;
wire            n2603;
wire            n2604;
wire            n2605;
wire            n2606;
wire            n2607;
wire            n2608;
wire            n2609;
wire            n261;
wire            n2610;
wire            n2611;
wire            n2612;
wire            n2613;
wire            n2614;
wire            n2615;
wire            n2616;
wire            n2617;
wire            n2618;
wire            n2619;
wire      [7:0] n262;
wire            n2620;
wire            n2621;
wire            n2622;
wire            n2623;
wire            n2624;
wire            n2625;
wire            n2626;
wire            n2627;
wire            n2628;
wire            n2629;
wire            n263;
wire            n2630;
wire            n2631;
wire            n2632;
wire            n2633;
wire            n2634;
wire            n2635;
wire            n2636;
wire            n2637;
wire            n2638;
wire            n2639;
wire            n264;
wire            n2640;
wire            n2641;
wire            n2642;
wire            n2643;
wire            n2644;
wire            n2645;
wire            n2646;
wire            n2647;
wire            n2648;
wire            n2649;
wire            n265;
wire            n2650;
wire            n2651;
wire            n2652;
wire            n2653;
wire            n2654;
wire            n2655;
wire            n2656;
wire            n2657;
wire            n2658;
wire            n2659;
wire            n266;
wire            n2660;
wire            n2661;
wire            n2662;
wire            n2663;
wire            n2664;
wire            n2665;
wire            n2666;
wire            n2667;
wire            n2668;
wire            n2669;
wire            n267;
wire            n2670;
wire            n2671;
wire            n2672;
wire            n2673;
wire            n2674;
wire            n2675;
wire            n2676;
wire            n2677;
wire            n2678;
wire            n2679;
wire            n268;
wire            n2680;
wire            n2681;
wire            n2682;
wire            n2683;
wire            n2684;
wire            n2685;
wire            n2686;
wire            n2687;
wire            n2688;
wire            n2689;
wire            n269;
wire            n2690;
wire            n2691;
wire            n2692;
wire            n2693;
wire            n2694;
wire            n2695;
wire            n2696;
wire            n2697;
wire            n2698;
wire            n2699;
wire            n27;
wire            n270;
wire            n2700;
wire            n2701;
wire            n2702;
wire            n2703;
wire            n2704;
wire            n2705;
wire            n2706;
wire            n2707;
wire            n2708;
wire            n2709;
wire            n271;
wire            n2710;
wire            n2711;
wire            n2712;
wire            n2713;
wire            n2714;
wire            n2715;
wire            n2716;
wire            n2717;
wire            n2718;
wire            n2719;
wire            n272;
wire            n2720;
wire            n2721;
wire            n2722;
wire            n2723;
wire            n2724;
wire            n2725;
wire            n2726;
wire            n2727;
wire            n2728;
wire            n2729;
wire            n273;
wire            n2730;
wire            n2731;
wire            n2732;
wire            n2733;
wire            n2734;
wire            n2735;
wire            n2736;
wire            n2737;
wire            n2738;
wire            n2739;
wire            n274;
wire            n2740;
wire            n2741;
wire            n2742;
wire            n2743;
wire            n2744;
wire            n2745;
wire            n2746;
wire            n2747;
wire            n2748;
wire            n2749;
wire            n275;
wire            n2750;
wire            n2751;
wire            n2752;
wire            n2753;
wire            n2754;
wire            n2755;
wire            n2756;
wire            n2757;
wire            n2758;
wire            n2759;
wire            n276;
wire            n2760;
wire            n2761;
wire            n2762;
wire            n2763;
wire            n2764;
wire            n2765;
wire            n2766;
wire            n2767;
wire            n2768;
wire            n2769;
wire            n277;
wire            n2770;
wire            n2771;
wire            n2772;
wire            n2773;
wire            n2774;
wire            n2775;
wire            n2776;
wire            n2777;
wire            n2778;
wire            n2779;
wire            n278;
wire            n2780;
wire            n2781;
wire            n2782;
wire            n2783;
wire            n2784;
wire            n2785;
wire            n2786;
wire            n2787;
wire            n2788;
wire            n2789;
wire            n279;
wire            n2790;
wire            n2791;
wire            n2792;
wire            n2793;
wire            n2794;
wire            n2795;
wire            n2796;
wire            n2797;
wire            n2798;
wire            n2799;
wire            n28;
wire            n280;
wire            n2800;
wire            n2801;
wire            n2802;
wire            n2803;
wire            n2804;
wire            n2805;
wire            n2806;
wire            n2807;
wire            n2808;
wire            n2809;
wire            n281;
wire            n2810;
wire            n2811;
wire            n2812;
wire            n2813;
wire            n2814;
wire            n2815;
wire            n2816;
wire            n2817;
wire            n2818;
wire            n2819;
wire            n282;
wire            n2820;
wire            n2821;
wire            n2822;
wire            n2823;
wire            n2824;
wire            n2825;
wire            n2826;
wire            n2827;
wire            n2828;
wire            n2829;
wire            n283;
wire            n2830;
wire            n2831;
wire            n2832;
wire            n2833;
wire            n2834;
wire            n2835;
wire            n2836;
wire            n2837;
wire            n2838;
wire            n2839;
wire      [7:0] n284;
wire            n2840;
wire            n2841;
wire            n2842;
wire            n2843;
wire            n2844;
wire            n2845;
wire            n2846;
wire            n2847;
wire            n2848;
wire            n2849;
wire            n285;
wire            n2850;
wire            n2851;
wire            n2852;
wire            n2853;
wire            n2854;
wire            n2855;
wire            n2856;
wire            n2857;
wire            n2858;
wire            n2859;
wire            n286;
wire            n2860;
wire            n2861;
wire            n2862;
wire            n2863;
wire            n2864;
wire            n2865;
wire            n2866;
wire            n2867;
wire            n2868;
wire            n2869;
wire            n287;
wire            n2870;
wire            n2871;
wire            n2872;
wire            n2873;
wire            n2874;
wire            n2875;
wire            n2876;
wire            n2877;
wire            n2878;
wire            n2879;
wire            n288;
wire            n2880;
wire            n2881;
wire            n2882;
wire            n2883;
wire            n2884;
wire            n2885;
wire            n2886;
wire            n2887;
wire            n2888;
wire            n2889;
wire            n289;
wire            n2890;
wire            n2891;
wire            n2892;
wire            n2893;
wire            n2894;
wire            n2895;
wire            n2896;
wire            n2897;
wire            n2898;
wire            n2899;
wire            n29;
wire            n290;
wire            n2900;
wire            n2901;
wire            n2902;
wire            n2903;
wire            n2904;
wire            n2905;
wire            n2906;
wire            n2907;
wire            n2908;
wire            n2909;
wire            n291;
wire            n2910;
wire            n2911;
wire            n2912;
wire            n2913;
wire            n2914;
wire            n2915;
wire            n2916;
wire            n2917;
wire            n2918;
wire            n2919;
wire            n292;
wire            n2920;
wire            n2921;
wire            n2922;
wire            n2923;
wire            n2924;
wire            n2925;
wire            n2926;
wire            n2927;
wire            n2928;
wire            n2929;
wire            n293;
wire            n2930;
wire            n2931;
wire            n2932;
wire            n2933;
wire            n2934;
wire            n2935;
wire            n2936;
wire            n2937;
wire            n2938;
wire            n2939;
wire            n294;
wire            n2940;
wire            n2941;
wire            n2942;
wire            n2943;
wire            n2944;
wire            n2945;
wire            n2946;
wire            n2947;
wire            n2948;
wire            n2949;
wire            n295;
wire            n2950;
wire            n2951;
wire            n2952;
wire            n2953;
wire            n2954;
wire            n2955;
wire            n2956;
wire            n2957;
wire            n2958;
wire            n2959;
wire            n296;
wire            n2960;
wire            n2961;
wire            n2962;
wire            n2963;
wire            n2964;
wire            n2965;
wire            n2966;
wire            n2967;
wire            n2968;
wire            n2969;
wire            n297;
wire            n2970;
wire            n2971;
wire            n2972;
wire            n2973;
wire            n2974;
wire            n2975;
wire            n2976;
wire            n2977;
wire            n2978;
wire            n2979;
wire            n298;
wire            n2980;
wire            n2981;
wire            n2982;
wire            n2983;
wire            n2984;
wire            n2985;
wire            n2986;
wire            n2987;
wire            n2988;
wire            n2989;
wire            n299;
wire            n2990;
wire            n2991;
wire            n2992;
wire            n2993;
wire            n2994;
wire            n2995;
wire            n2996;
wire            n2997;
wire            n2998;
wire            n2999;
wire            n3;
wire            n30;
wire            n300;
wire            n3000;
wire            n3001;
wire            n3002;
wire            n3003;
wire            n3004;
wire            n3005;
wire            n3006;
wire            n3007;
wire            n3008;
wire            n3009;
wire            n301;
wire            n3010;
wire            n3011;
wire            n3012;
wire            n3013;
wire            n3014;
wire            n3015;
wire            n3016;
wire            n3017;
wire            n3018;
wire            n3019;
wire            n302;
wire            n3020;
wire            n3021;
wire            n3022;
wire            n3023;
wire            n3024;
wire            n3025;
wire            n3026;
wire            n3027;
wire            n3028;
wire            n3029;
wire            n303;
wire            n3030;
wire            n3031;
wire            n3032;
wire            n3033;
wire            n3034;
wire            n3035;
wire            n3036;
wire            n3037;
wire            n3038;
wire            n3039;
wire            n304;
wire            n3040;
wire            n3041;
wire            n3042;
wire            n3043;
wire            n3044;
wire            n3045;
wire            n3046;
wire            n3047;
wire            n3048;
wire            n3049;
wire            n305;
wire            n3050;
wire            n3051;
wire            n3052;
wire            n3053;
wire            n3054;
wire            n3055;
wire            n3056;
wire            n3057;
wire            n3058;
wire            n3059;
wire      [7:0] n306;
wire            n3060;
wire            n3061;
wire            n3062;
wire            n3063;
wire            n3064;
wire            n3065;
wire            n3066;
wire            n3067;
wire            n3068;
wire            n3069;
wire            n307;
wire            n3070;
wire            n3071;
wire            n3072;
wire            n3073;
wire            n3074;
wire            n3075;
wire            n3076;
wire            n3077;
wire            n3078;
wire            n3079;
wire            n308;
wire            n3080;
wire            n3081;
wire            n3082;
wire            n3083;
wire            n3084;
wire            n3085;
wire            n3086;
wire            n3087;
wire            n3088;
wire            n3089;
wire            n309;
wire            n3090;
wire            n3091;
wire            n3092;
wire            n3093;
wire            n3094;
wire            n3095;
wire            n3096;
wire            n3097;
wire            n3098;
wire            n3099;
wire            n31;
wire            n310;
wire            n3100;
wire            n3101;
wire            n3102;
wire            n3103;
wire            n3104;
wire            n3105;
wire            n3106;
wire            n3107;
wire            n3108;
wire            n3109;
wire            n311;
wire            n3110;
wire            n3111;
wire            n3112;
wire            n3113;
wire            n3114;
wire            n3115;
wire            n3116;
wire            n3117;
wire            n3118;
wire            n3119;
wire            n312;
wire            n3120;
wire            n3121;
wire            n3122;
wire            n3123;
wire            n3124;
wire            n3125;
wire            n3126;
wire            n3127;
wire            n3128;
wire            n3129;
wire            n313;
wire            n3130;
wire            n3131;
wire            n3132;
wire            n3133;
wire            n3134;
wire            n3135;
wire            n3136;
wire            n3137;
wire            n3138;
wire            n3139;
wire            n314;
wire            n3140;
wire            n3141;
wire            n3142;
wire            n3143;
wire            n3144;
wire            n3145;
wire            n3146;
wire            n3147;
wire            n3148;
wire            n3149;
wire            n315;
wire            n3150;
wire            n3151;
wire            n3152;
wire            n3153;
wire            n3154;
wire            n3155;
wire            n3156;
wire            n3157;
wire            n3158;
wire            n3159;
wire            n316;
wire            n3160;
wire            n3161;
wire            n3162;
wire            n3163;
wire            n3164;
wire            n3165;
wire            n3166;
wire            n3167;
wire            n3168;
wire            n3169;
wire            n317;
wire            n3170;
wire            n3171;
wire            n3172;
wire            n3173;
wire            n3174;
wire            n3175;
wire            n3176;
wire            n3177;
wire            n3178;
wire            n3179;
wire            n318;
wire            n3180;
wire            n3181;
wire            n3182;
wire            n3183;
wire            n3184;
wire            n3185;
wire            n3186;
wire            n3187;
wire            n3188;
wire            n3189;
wire            n319;
wire            n3190;
wire            n3191;
wire            n3192;
wire            n3193;
wire            n3194;
wire            n3195;
wire            n3196;
wire            n3197;
wire            n3198;
wire            n3199;
wire            n32;
wire            n320;
wire            n3200;
wire            n3201;
wire            n3202;
wire            n3203;
wire            n3204;
wire            n3205;
wire            n3206;
wire            n3207;
wire            n3208;
wire            n3209;
wire            n321;
wire            n3210;
wire            n3211;
wire            n3212;
wire            n3213;
wire            n3214;
wire            n3215;
wire            n3216;
wire            n3217;
wire            n3218;
wire            n3219;
wire            n322;
wire            n3220;
wire            n3221;
wire            n3222;
wire            n3223;
wire            n3224;
wire            n3225;
wire            n3226;
wire            n3227;
wire            n3228;
wire            n3229;
wire            n323;
wire            n3230;
wire            n3231;
wire            n3232;
wire            n3233;
wire            n3234;
wire            n3235;
wire            n3236;
wire            n3237;
wire            n3238;
wire            n3239;
wire            n324;
wire            n3240;
wire            n3241;
wire            n3242;
wire            n3243;
wire            n3244;
wire            n3245;
wire            n3246;
wire            n3247;
wire            n3248;
wire            n3249;
wire            n325;
wire            n3250;
wire            n3251;
wire            n3252;
wire            n3253;
wire            n3254;
wire            n3255;
wire            n3256;
wire            n3257;
wire            n3258;
wire            n3259;
wire            n326;
wire            n3260;
wire            n3261;
wire            n3262;
wire            n3263;
wire            n3264;
wire            n3265;
wire            n3266;
wire            n3267;
wire            n3268;
wire            n3269;
wire            n327;
wire            n3270;
wire            n3271;
wire            n3272;
wire            n3273;
wire            n3274;
wire            n3275;
wire            n3276;
wire            n3277;
wire            n3278;
wire            n3279;
wire      [7:0] n328;
wire            n3280;
wire            n3281;
wire            n3282;
wire            n3283;
wire            n3284;
wire            n3285;
wire            n3286;
wire            n3287;
wire            n3288;
wire            n3289;
wire            n329;
wire            n3290;
wire            n3291;
wire            n3292;
wire            n3293;
wire            n3294;
wire            n3295;
wire            n3296;
wire            n3297;
wire            n3298;
wire            n3299;
wire            n33;
wire            n330;
wire            n3300;
wire            n3301;
wire            n3302;
wire            n3303;
wire            n3304;
wire            n3305;
wire            n3306;
wire            n3307;
wire            n3308;
wire            n3309;
wire            n331;
wire            n3310;
wire            n3311;
wire            n3312;
wire            n3313;
wire            n3314;
wire            n3315;
wire            n3316;
wire            n3317;
wire            n3318;
wire            n3319;
wire            n332;
wire            n3320;
wire            n3321;
wire            n3322;
wire            n3323;
wire            n3324;
wire            n3325;
wire            n3326;
wire            n3327;
wire            n3328;
wire            n3329;
wire            n333;
wire            n3330;
wire            n3331;
wire            n3332;
wire            n3333;
wire            n3334;
wire            n3335;
wire            n3336;
wire            n3337;
wire            n3338;
wire            n3339;
wire            n334;
wire            n3340;
wire            n3341;
wire            n3342;
wire            n3343;
wire            n3344;
wire            n3345;
wire            n3346;
wire            n3347;
wire            n3348;
wire            n3349;
wire            n335;
wire            n3350;
wire            n3351;
wire            n3352;
wire            n3353;
wire            n3354;
wire            n3355;
wire            n3356;
wire            n3357;
wire            n3358;
wire            n3359;
wire            n336;
wire            n3360;
wire            n3361;
wire            n3362;
wire            n3363;
wire            n3364;
wire            n3365;
wire            n3366;
wire            n3367;
wire            n3368;
wire            n3369;
wire            n337;
wire            n3370;
wire            n3371;
wire            n3372;
wire            n3373;
wire            n3374;
wire            n3375;
wire            n3376;
wire            n3377;
wire            n3378;
wire            n3379;
wire            n338;
wire            n3380;
wire            n3381;
wire            n3382;
wire            n3383;
wire            n3384;
wire            n3385;
wire            n3386;
wire            n3387;
wire            n3388;
wire            n3389;
wire            n339;
wire            n3390;
wire            n3391;
wire            n3392;
wire            n3393;
wire            n3394;
wire            n3395;
wire            n3396;
wire            n3397;
wire            n3398;
wire            n3399;
wire            n34;
wire            n340;
wire            n3400;
wire            n3401;
wire            n3402;
wire            n3403;
wire            n3404;
wire            n3405;
wire            n3406;
wire            n3407;
wire            n3408;
wire            n3409;
wire            n341;
wire            n3410;
wire            n3411;
wire            n3412;
wire            n3413;
wire            n3414;
wire            n3415;
wire            n3416;
wire            n3417;
wire            n3418;
wire            n3419;
wire            n342;
wire            n3420;
wire            n3421;
wire            n3422;
wire            n3423;
wire            n3424;
wire            n3425;
wire            n3426;
wire            n3427;
wire            n3428;
wire            n3429;
wire            n343;
wire            n3430;
wire            n3431;
wire            n3432;
wire            n3433;
wire            n3434;
wire            n3435;
wire            n3436;
wire            n3437;
wire            n3438;
wire            n3439;
wire            n344;
wire            n3440;
wire            n3441;
wire            n3442;
wire            n3443;
wire            n3444;
wire            n3445;
wire            n3446;
wire            n3447;
wire            n3448;
wire            n3449;
wire            n345;
wire            n3450;
wire            n3451;
wire            n3452;
wire            n3453;
wire            n3454;
wire            n3455;
wire            n3456;
wire            n3457;
wire            n3458;
wire            n3459;
wire            n346;
wire            n3460;
wire            n3461;
wire            n3462;
wire            n3463;
wire            n3464;
wire            n3465;
wire            n3466;
wire            n3467;
wire            n3468;
wire            n3469;
wire            n347;
wire            n3470;
wire            n3471;
wire            n3472;
wire            n3473;
wire            n3474;
wire            n3475;
wire            n3476;
wire            n3477;
wire            n3478;
wire            n3479;
wire            n348;
wire            n3480;
wire            n3481;
wire            n3482;
wire            n3483;
wire            n3484;
wire            n3485;
wire            n3486;
wire            n3487;
wire            n3488;
wire            n3489;
wire            n349;
wire            n3490;
wire            n3491;
wire            n3492;
wire            n3493;
wire            n3494;
wire            n35;
wire            n350;
wire      [7:0] n351;
wire            n352;
wire            n353;
wire            n354;
wire            n355;
wire            n356;
wire            n357;
wire            n358;
wire            n359;
wire            n36;
wire            n360;
wire            n361;
wire            n362;
wire            n363;
wire            n364;
wire            n365;
wire            n366;
wire            n367;
wire            n368;
wire            n369;
wire            n37;
wire            n370;
wire            n371;
wire            n372;
wire            n373;
wire            n374;
wire            n375;
wire            n376;
wire            n377;
wire            n378;
wire            n379;
wire            n38;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n39;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n4;
wire            n40;
wire            n400;
wire            n401;
wire            n402;
wire            n403;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n41;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n42;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n43;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n44;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire            n447;
wire            n448;
wire            n449;
wire            n45;
wire            n450;
wire            n451;
wire            n452;
wire            n453;
wire            n454;
wire            n455;
wire            n456;
wire            n457;
wire            n458;
wire            n459;
wire            n46;
wire            n460;
wire            n461;
wire            n462;
wire            n463;
wire            n464;
wire            n465;
wire            n466;
wire            n467;
wire            n468;
wire            n469;
wire            n47;
wire            n470;
wire            n471;
wire            n472;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire            n478;
wire            n479;
wire            n48;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n49;
wire            n490;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n5;
wire            n50;
wire            n500;
wire            n501;
wire            n502;
wire            n503;
wire            n504;
wire            n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n51;
wire            n510;
wire            n511;
wire            n512;
wire            n513;
wire            n514;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
wire            n519;
wire            n52;
wire            n520;
wire            n521;
wire            n522;
wire            n523;
wire            n524;
wire            n525;
wire            n526;
wire            n527;
wire            n528;
wire            n529;
wire            n53;
wire            n530;
wire            n531;
wire            n532;
wire            n533;
wire            n534;
wire            n535;
wire            n536;
wire            n537;
wire            n538;
wire            n539;
wire            n54;
wire            n540;
wire            n541;
wire            n542;
wire            n543;
wire            n544;
wire            n545;
wire            n546;
wire            n547;
wire            n548;
wire            n549;
wire            n55;
wire            n550;
wire            n551;
wire            n552;
wire            n553;
wire            n554;
wire            n555;
wire            n556;
wire            n557;
wire            n558;
wire            n559;
wire            n56;
wire            n560;
wire            n561;
wire            n562;
wire            n563;
wire            n564;
wire            n565;
wire            n566;
wire            n567;
wire            n568;
wire            n569;
wire            n57;
wire            n570;
wire            n571;
wire            n572;
wire            n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n58;
wire            n580;
wire            n581;
wire            n582;
wire            n583;
wire            n584;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n589;
wire            n59;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n6;
wire            n60;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n61;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n62;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n63;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n64;
wire            n640;
wire            n641;
wire      [7:0] n642;
wire      [7:0] n643;
wire      [7:0] n644;
wire      [7:0] n645;
wire      [7:0] n646;
wire      [7:0] n647;
wire      [7:0] n648;
wire      [7:0] n649;
wire            n65;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire            n658;
wire            n659;
wire            n66;
wire            n660;
wire            n661;
wire            n662;
wire            n663;
wire            n664;
wire            n665;
wire            n666;
wire            n667;
wire            n668;
wire            n669;
wire            n67;
wire            n670;
wire            n671;
wire            n672;
wire            n673;
wire            n674;
wire            n675;
wire            n676;
wire            n677;
wire            n678;
wire            n679;
wire            n68;
wire            n680;
wire            n681;
wire            n682;
wire            n683;
wire            n684;
wire            n685;
wire            n686;
wire            n687;
wire            n688;
wire            n689;
wire            n69;
wire            n690;
wire            n691;
wire            n692;
wire            n693;
wire            n694;
wire            n695;
wire            n696;
wire            n697;
wire            n698;
wire            n699;
wire            n7;
wire            n70;
wire            n700;
wire            n701;
wire            n702;
wire            n703;
wire            n704;
wire            n705;
wire            n706;
wire            n707;
wire            n708;
wire            n709;
wire            n71;
wire            n710;
wire            n711;
wire            n712;
wire            n713;
wire            n714;
wire            n715;
wire            n716;
wire            n717;
wire            n718;
wire            n719;
wire            n72;
wire            n720;
wire            n721;
wire            n722;
wire            n723;
wire            n724;
wire            n725;
wire            n726;
wire            n727;
wire            n728;
wire            n729;
wire            n73;
wire            n730;
wire            n731;
wire            n732;
wire     [15:0] n733;
wire     [15:0] n734;
wire            n735;
wire     [15:0] n736;
wire            n737;
wire            n738;
wire            n739;
wire            n74;
wire            n740;
wire            n741;
wire            n742;
wire            n743;
wire            n744;
wire            n745;
wire            n746;
wire            n747;
wire            n748;
wire            n749;
wire            n75;
wire            n750;
wire            n751;
wire            n752;
wire            n753;
wire            n754;
wire            n755;
wire            n756;
wire            n757;
wire            n758;
wire            n759;
wire            n76;
wire            n760;
wire            n761;
wire            n762;
wire            n763;
wire            n764;
wire            n765;
wire            n766;
wire            n767;
wire            n768;
wire            n769;
wire            n77;
wire            n770;
wire            n771;
wire            n772;
wire            n773;
wire            n774;
wire            n775;
wire            n776;
wire            n777;
wire            n778;
wire            n779;
wire            n78;
wire            n780;
wire            n781;
wire            n782;
wire            n783;
wire            n784;
wire            n785;
wire            n786;
wire            n787;
wire            n788;
wire            n789;
wire            n79;
wire            n790;
wire            n791;
wire            n792;
wire            n793;
wire            n794;
wire            n795;
wire            n796;
wire            n797;
wire            n798;
wire            n799;
wire            n8;
wire            n80;
wire            n800;
wire            n801;
wire            n802;
wire            n803;
wire            n804;
wire            n805;
wire            n806;
wire            n807;
wire            n808;
wire            n809;
wire            n81;
wire            n810;
wire            n811;
wire            n812;
wire            n813;
wire            n814;
wire            n815;
wire            n816;
wire            n817;
wire            n818;
wire            n819;
wire            n82;
wire            n820;
wire    [159:0] n821;
wire    [159:0] n823;
wire    [159:0] n824;
wire      [7:0] n825;
wire     [15:0] n826;
wire      [7:0] n827;
wire     [15:0] n828;
wire            n829;
wire            n83;
wire            n830;
wire            n831;
wire            n832;
wire            n833;
wire            n834;
wire            n835;
wire            n836;
wire            n837;
wire            n838;
wire            n839;
wire            n84;
wire            n840;
wire            n841;
wire            n842;
wire            n843;
wire            n844;
wire            n845;
wire            n846;
wire            n847;
wire            n848;
wire            n849;
wire            n85;
wire            n850;
wire            n851;
wire            n852;
wire            n853;
wire            n854;
wire            n855;
wire            n856;
wire            n857;
wire            n858;
wire            n859;
wire            n86;
wire            n860;
wire            n861;
wire            n862;
wire            n863;
wire            n864;
wire            n865;
wire            n866;
wire            n867;
wire            n868;
wire            n869;
wire            n87;
wire            n870;
wire            n871;
wire            n872;
wire            n873;
wire            n874;
wire            n875;
wire            n876;
wire            n877;
wire            n878;
wire            n879;
wire            n88;
wire            n880;
wire            n881;
wire            n882;
wire            n883;
wire            n884;
wire            n885;
wire            n886;
wire            n887;
wire            n888;
wire            n889;
wire            n89;
wire            n890;
wire            n891;
wire            n892;
wire            n893;
wire            n894;
wire            n895;
wire            n896;
wire            n897;
wire            n898;
wire            n899;
wire            n9;
wire            n90;
wire            n900;
wire            n901;
wire            n902;
wire            n903;
wire            n904;
wire            n905;
wire            n906;
wire            n907;
wire            n908;
wire            n909;
wire            n91;
wire            n910;
wire            n911;
wire     [15:0] n912;
wire     [15:0] n913;
wire      [7:0] n916;
wire     [15:0] n917;
wire            n92;
wire      [7:0] n920;
wire     [15:0] n921;
wire     [15:0] n922;
wire      [7:0] n925;
wire     [23:0] n926;
wire     [15:0] n927;
wire            n93;
wire      [7:0] n930;
wire     [31:0] n931;
wire     [15:0] n932;
wire      [7:0] n935;
wire     [39:0] n936;
wire     [15:0] n937;
wire            n94;
wire      [7:0] n940;
wire     [47:0] n941;
wire     [15:0] n942;
wire      [7:0] n945;
wire     [55:0] n946;
wire     [15:0] n947;
wire            n95;
wire      [7:0] n950;
wire     [63:0] n951;
wire     [15:0] n952;
wire      [7:0] n955;
wire     [71:0] n956;
wire     [15:0] n957;
wire            n96;
wire      [7:0] n960;
wire     [79:0] n961;
wire     [15:0] n962;
wire      [7:0] n965;
wire     [87:0] n966;
wire     [15:0] n967;
wire            n97;
wire      [7:0] n970;
wire     [95:0] n971;
wire     [15:0] n972;
wire      [7:0] n975;
wire    [103:0] n976;
wire     [15:0] n977;
wire            n98;
wire      [7:0] n980;
wire    [111:0] n981;
wire     [15:0] n982;
wire      [7:0] n985;
wire    [119:0] n986;
wire     [15:0] n987;
wire            n99;
wire      [7:0] n990;
wire    [127:0] n991;
wire     [15:0] n992;
wire      [7:0] n995;
wire    [135:0] n996;
wire     [15:0] n997;
wire            rst;
assign __ILA_sha_valid__ = 1'b1 ;
assign n0 =  ( sha_state ) == ( 3'd0 )  ;
assign n1 =  ( cmd ) == ( 2'd1 )  ;
assign n2 =  ( n0 ) & (n1 )  ;
assign n3 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n4 =  ( n2 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__0__ = n4 ;
assign __ILA_sha_acc_decode__[0] = __ILA_sha_decode_of_I__DOT__0__ ;
assign n5 =  ( sha_state ) == ( 3'd1 )  ;
assign n6 =  ( n5 ) & (n1 )  ;
assign n7 =  ( n6 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__1__ = n7 ;
assign __ILA_sha_acc_decode__[1] = __ILA_sha_decode_of_I__DOT__1__ ;
assign n8 =  ( sha_state ) == ( 3'd2 )  ;
assign n9 =  ( n8 ) & (n1 )  ;
assign n10 =  ( n9 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__2__ = n10 ;
assign __ILA_sha_acc_decode__[2] = __ILA_sha_decode_of_I__DOT__2__ ;
assign n11 =  ( sha_state ) == ( 3'd3 )  ;
assign n12 =  ( n11 ) & (n1 )  ;
assign n13 =  ( n12 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__3__ = n13 ;
assign __ILA_sha_acc_decode__[3] = __ILA_sha_decode_of_I__DOT__3__ ;
assign n14 =  ( sha_state ) == ( 3'd4 )  ;
assign n15 =  ( n14 ) & (n1 )  ;
assign n16 =  ( n15 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__4__ = n16 ;
assign __ILA_sha_acc_decode__[4] = __ILA_sha_decode_of_I__DOT__4__ ;
assign n17 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n18 =  ( n2 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__5__ = n18 ;
assign __ILA_sha_acc_decode__[5] = __ILA_sha_decode_of_I__DOT__5__ ;
assign n19 =  ( n6 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__6__ = n19 ;
assign __ILA_sha_acc_decode__[6] = __ILA_sha_decode_of_I__DOT__6__ ;
assign n20 =  ( n9 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__7__ = n20 ;
assign __ILA_sha_acc_decode__[7] = __ILA_sha_decode_of_I__DOT__7__ ;
assign n21 =  ( n12 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__8__ = n21 ;
assign __ILA_sha_acc_decode__[8] = __ILA_sha_decode_of_I__DOT__8__ ;
assign n22 =  ( n15 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__9__ = n22 ;
assign __ILA_sha_acc_decode__[9] = __ILA_sha_decode_of_I__DOT__9__ ;
assign n23 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n24 =  ( n2 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__10__ = n24 ;
assign __ILA_sha_acc_decode__[10] = __ILA_sha_decode_of_I__DOT__10__ ;
assign n25 =  ( n6 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__11__ = n25 ;
assign __ILA_sha_acc_decode__[11] = __ILA_sha_decode_of_I__DOT__11__ ;
assign n26 =  ( n9 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__12__ = n26 ;
assign __ILA_sha_acc_decode__[12] = __ILA_sha_decode_of_I__DOT__12__ ;
assign n27 =  ( n12 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__13__ = n27 ;
assign __ILA_sha_acc_decode__[13] = __ILA_sha_decode_of_I__DOT__13__ ;
assign n28 =  ( n15 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__14__ = n28 ;
assign __ILA_sha_acc_decode__[14] = __ILA_sha_decode_of_I__DOT__14__ ;
assign n29 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n30 =  ( n2 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__15__ = n30 ;
assign __ILA_sha_acc_decode__[15] = __ILA_sha_decode_of_I__DOT__15__ ;
assign n31 =  ( n6 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__16__ = n31 ;
assign __ILA_sha_acc_decode__[16] = __ILA_sha_decode_of_I__DOT__16__ ;
assign n32 =  ( n9 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__17__ = n32 ;
assign __ILA_sha_acc_decode__[17] = __ILA_sha_decode_of_I__DOT__17__ ;
assign n33 =  ( n12 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__18__ = n33 ;
assign __ILA_sha_acc_decode__[18] = __ILA_sha_decode_of_I__DOT__18__ ;
assign n34 =  ( n15 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__19__ = n34 ;
assign __ILA_sha_acc_decode__[19] = __ILA_sha_decode_of_I__DOT__19__ ;
assign n35 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n36 =  ( n2 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__20__ = n36 ;
assign __ILA_sha_acc_decode__[20] = __ILA_sha_decode_of_I__DOT__20__ ;
assign n37 =  ( n6 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__21__ = n37 ;
assign __ILA_sha_acc_decode__[21] = __ILA_sha_decode_of_I__DOT__21__ ;
assign n38 =  ( n9 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__22__ = n38 ;
assign __ILA_sha_acc_decode__[22] = __ILA_sha_decode_of_I__DOT__22__ ;
assign n39 =  ( n12 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__23__ = n39 ;
assign __ILA_sha_acc_decode__[23] = __ILA_sha_decode_of_I__DOT__23__ ;
assign n40 =  ( n15 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__24__ = n40 ;
assign __ILA_sha_acc_decode__[24] = __ILA_sha_decode_of_I__DOT__24__ ;
assign n41 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n42 =  ( n2 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__25__ = n42 ;
assign __ILA_sha_acc_decode__[25] = __ILA_sha_decode_of_I__DOT__25__ ;
assign n43 =  ( n6 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__26__ = n43 ;
assign __ILA_sha_acc_decode__[26] = __ILA_sha_decode_of_I__DOT__26__ ;
assign n44 =  ( n9 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__27__ = n44 ;
assign __ILA_sha_acc_decode__[27] = __ILA_sha_decode_of_I__DOT__27__ ;
assign n45 =  ( n12 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__28__ = n45 ;
assign __ILA_sha_acc_decode__[28] = __ILA_sha_decode_of_I__DOT__28__ ;
assign n46 =  ( n15 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__29__ = n46 ;
assign __ILA_sha_acc_decode__[29] = __ILA_sha_decode_of_I__DOT__29__ ;
assign n47 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n48 =  ( n2 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__30__ = n48 ;
assign __ILA_sha_acc_decode__[30] = __ILA_sha_decode_of_I__DOT__30__ ;
assign n49 =  ( n6 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__31__ = n49 ;
assign __ILA_sha_acc_decode__[31] = __ILA_sha_decode_of_I__DOT__31__ ;
assign n50 =  ( n9 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__32__ = n50 ;
assign __ILA_sha_acc_decode__[32] = __ILA_sha_decode_of_I__DOT__32__ ;
assign n51 =  ( n12 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__33__ = n51 ;
assign __ILA_sha_acc_decode__[33] = __ILA_sha_decode_of_I__DOT__33__ ;
assign n52 =  ( n15 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__34__ = n52 ;
assign __ILA_sha_acc_decode__[34] = __ILA_sha_decode_of_I__DOT__34__ ;
assign n53 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n54 =  ( n2 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__35__ = n54 ;
assign __ILA_sha_acc_decode__[35] = __ILA_sha_decode_of_I__DOT__35__ ;
assign n55 =  ( n6 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__36__ = n55 ;
assign __ILA_sha_acc_decode__[36] = __ILA_sha_decode_of_I__DOT__36__ ;
assign n56 =  ( n9 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__37__ = n56 ;
assign __ILA_sha_acc_decode__[37] = __ILA_sha_decode_of_I__DOT__37__ ;
assign n57 =  ( n12 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__38__ = n57 ;
assign __ILA_sha_acc_decode__[38] = __ILA_sha_decode_of_I__DOT__38__ ;
assign n58 =  ( n15 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__39__ = n58 ;
assign __ILA_sha_acc_decode__[39] = __ILA_sha_decode_of_I__DOT__39__ ;
assign n59 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n60 =  ( n2 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__40__ = n60 ;
assign __ILA_sha_acc_decode__[40] = __ILA_sha_decode_of_I__DOT__40__ ;
assign n61 =  ( n6 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__41__ = n61 ;
assign __ILA_sha_acc_decode__[41] = __ILA_sha_decode_of_I__DOT__41__ ;
assign n62 =  ( n9 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__42__ = n62 ;
assign __ILA_sha_acc_decode__[42] = __ILA_sha_decode_of_I__DOT__42__ ;
assign n63 =  ( n12 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__43__ = n63 ;
assign __ILA_sha_acc_decode__[43] = __ILA_sha_decode_of_I__DOT__43__ ;
assign n64 =  ( n15 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__44__ = n64 ;
assign __ILA_sha_acc_decode__[44] = __ILA_sha_decode_of_I__DOT__44__ ;
assign n65 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n66 =  ( n2 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__45__ = n66 ;
assign __ILA_sha_acc_decode__[45] = __ILA_sha_decode_of_I__DOT__45__ ;
assign n67 =  ( n6 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__46__ = n67 ;
assign __ILA_sha_acc_decode__[46] = __ILA_sha_decode_of_I__DOT__46__ ;
assign n68 =  ( n9 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__47__ = n68 ;
assign __ILA_sha_acc_decode__[47] = __ILA_sha_decode_of_I__DOT__47__ ;
assign n69 =  ( n12 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__48__ = n69 ;
assign __ILA_sha_acc_decode__[48] = __ILA_sha_decode_of_I__DOT__48__ ;
assign n70 =  ( n15 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__49__ = n70 ;
assign __ILA_sha_acc_decode__[49] = __ILA_sha_decode_of_I__DOT__49__ ;
assign n71 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n72 =  ( n2 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__50__ = n72 ;
assign __ILA_sha_acc_decode__[50] = __ILA_sha_decode_of_I__DOT__50__ ;
assign n73 =  ( n6 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__51__ = n73 ;
assign __ILA_sha_acc_decode__[51] = __ILA_sha_decode_of_I__DOT__51__ ;
assign n74 =  ( n9 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__52__ = n74 ;
assign __ILA_sha_acc_decode__[52] = __ILA_sha_decode_of_I__DOT__52__ ;
assign n75 =  ( n12 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__53__ = n75 ;
assign __ILA_sha_acc_decode__[53] = __ILA_sha_decode_of_I__DOT__53__ ;
assign n76 =  ( n15 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__54__ = n76 ;
assign __ILA_sha_acc_decode__[54] = __ILA_sha_decode_of_I__DOT__54__ ;
assign n77 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n78 =  ( n2 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__55__ = n78 ;
assign __ILA_sha_acc_decode__[55] = __ILA_sha_decode_of_I__DOT__55__ ;
assign n79 =  ( n6 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__56__ = n79 ;
assign __ILA_sha_acc_decode__[56] = __ILA_sha_decode_of_I__DOT__56__ ;
assign n80 =  ( n9 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__57__ = n80 ;
assign __ILA_sha_acc_decode__[57] = __ILA_sha_decode_of_I__DOT__57__ ;
assign n81 =  ( n12 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__58__ = n81 ;
assign __ILA_sha_acc_decode__[58] = __ILA_sha_decode_of_I__DOT__58__ ;
assign n82 =  ( n15 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__59__ = n82 ;
assign __ILA_sha_acc_decode__[59] = __ILA_sha_decode_of_I__DOT__59__ ;
assign n83 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n84 =  ( n2 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__60__ = n84 ;
assign __ILA_sha_acc_decode__[60] = __ILA_sha_decode_of_I__DOT__60__ ;
assign n85 =  ( n6 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__61__ = n85 ;
assign __ILA_sha_acc_decode__[61] = __ILA_sha_decode_of_I__DOT__61__ ;
assign n86 =  ( n9 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__62__ = n86 ;
assign __ILA_sha_acc_decode__[62] = __ILA_sha_decode_of_I__DOT__62__ ;
assign n87 =  ( n12 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__63__ = n87 ;
assign __ILA_sha_acc_decode__[63] = __ILA_sha_decode_of_I__DOT__63__ ;
assign n88 =  ( n15 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__64__ = n88 ;
assign __ILA_sha_acc_decode__[64] = __ILA_sha_decode_of_I__DOT__64__ ;
assign n89 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n90 =  ( n2 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__65__ = n90 ;
assign __ILA_sha_acc_decode__[65] = __ILA_sha_decode_of_I__DOT__65__ ;
assign n91 =  ( n6 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__66__ = n91 ;
assign __ILA_sha_acc_decode__[66] = __ILA_sha_decode_of_I__DOT__66__ ;
assign n92 =  ( n9 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__67__ = n92 ;
assign __ILA_sha_acc_decode__[67] = __ILA_sha_decode_of_I__DOT__67__ ;
assign n93 =  ( n12 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__68__ = n93 ;
assign __ILA_sha_acc_decode__[68] = __ILA_sha_decode_of_I__DOT__68__ ;
assign n94 =  ( n15 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__69__ = n94 ;
assign __ILA_sha_acc_decode__[69] = __ILA_sha_decode_of_I__DOT__69__ ;
assign n95 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n96 =  ( n2 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__70__ = n96 ;
assign __ILA_sha_acc_decode__[70] = __ILA_sha_decode_of_I__DOT__70__ ;
assign n97 =  ( n6 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__71__ = n97 ;
assign __ILA_sha_acc_decode__[71] = __ILA_sha_decode_of_I__DOT__71__ ;
assign n98 =  ( n9 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__72__ = n98 ;
assign __ILA_sha_acc_decode__[72] = __ILA_sha_decode_of_I__DOT__72__ ;
assign n99 =  ( n12 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__73__ = n99 ;
assign __ILA_sha_acc_decode__[73] = __ILA_sha_decode_of_I__DOT__73__ ;
assign n100 =  ( n15 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__74__ = n100 ;
assign __ILA_sha_acc_decode__[74] = __ILA_sha_decode_of_I__DOT__74__ ;
assign n101 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n102 =  ( n2 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__75__ = n102 ;
assign __ILA_sha_acc_decode__[75] = __ILA_sha_decode_of_I__DOT__75__ ;
assign n103 =  ( n6 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__76__ = n103 ;
assign __ILA_sha_acc_decode__[76] = __ILA_sha_decode_of_I__DOT__76__ ;
assign n104 =  ( n9 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__77__ = n104 ;
assign __ILA_sha_acc_decode__[77] = __ILA_sha_decode_of_I__DOT__77__ ;
assign n105 =  ( n12 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__78__ = n105 ;
assign __ILA_sha_acc_decode__[78] = __ILA_sha_decode_of_I__DOT__78__ ;
assign n106 =  ( n15 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__79__ = n106 ;
assign __ILA_sha_acc_decode__[79] = __ILA_sha_decode_of_I__DOT__79__ ;
assign n107 =  ( cmd ) == ( 2'd2 )  ;
assign n108 =  ( n0 ) & (n107 )  ;
assign n109 =  ( n108 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__80__ = n109 ;
assign __ILA_sha_acc_decode__[80] = __ILA_sha_decode_of_I__DOT__80__ ;
assign n110 =  ( n108 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__81__ = n110 ;
assign __ILA_sha_acc_decode__[81] = __ILA_sha_decode_of_I__DOT__81__ ;
assign n111 =  ( n108 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__82__ = n111 ;
assign __ILA_sha_acc_decode__[82] = __ILA_sha_decode_of_I__DOT__82__ ;
assign n112 =  ( n108 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__83__ = n112 ;
assign __ILA_sha_acc_decode__[83] = __ILA_sha_decode_of_I__DOT__83__ ;
assign n113 =  ( n108 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__84__ = n113 ;
assign __ILA_sha_acc_decode__[84] = __ILA_sha_decode_of_I__DOT__84__ ;
assign n114 =  ( n108 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__85__ = n114 ;
assign __ILA_sha_acc_decode__[85] = __ILA_sha_decode_of_I__DOT__85__ ;
assign n115 =  ( n108 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__86__ = n115 ;
assign __ILA_sha_acc_decode__[86] = __ILA_sha_decode_of_I__DOT__86__ ;
assign n116 =  ( n108 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__87__ = n116 ;
assign __ILA_sha_acc_decode__[87] = __ILA_sha_decode_of_I__DOT__87__ ;
assign n117 =  ( n108 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__88__ = n117 ;
assign __ILA_sha_acc_decode__[88] = __ILA_sha_decode_of_I__DOT__88__ ;
assign n118 =  ( n108 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__89__ = n118 ;
assign __ILA_sha_acc_decode__[89] = __ILA_sha_decode_of_I__DOT__89__ ;
assign n119 =  ( n108 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__90__ = n119 ;
assign __ILA_sha_acc_decode__[90] = __ILA_sha_decode_of_I__DOT__90__ ;
assign n120 =  ( n108 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__91__ = n120 ;
assign __ILA_sha_acc_decode__[91] = __ILA_sha_decode_of_I__DOT__91__ ;
assign n121 =  ( n108 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__92__ = n121 ;
assign __ILA_sha_acc_decode__[92] = __ILA_sha_decode_of_I__DOT__92__ ;
assign n122 =  ( n108 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__93__ = n122 ;
assign __ILA_sha_acc_decode__[93] = __ILA_sha_decode_of_I__DOT__93__ ;
assign n123 =  ( n108 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__94__ = n123 ;
assign __ILA_sha_acc_decode__[94] = __ILA_sha_decode_of_I__DOT__94__ ;
assign n124 =  ( n108 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__95__ = n124 ;
assign __ILA_sha_acc_decode__[95] = __ILA_sha_decode_of_I__DOT__95__ ;
assign n125 = ~ ( n1 )  ;
assign n126 =  ( n5 ) & (n125 )  ;
assign n127 =  ( n126 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__96__ = n127 ;
assign __ILA_sha_acc_decode__[96] = __ILA_sha_decode_of_I__DOT__96__ ;
assign n128 =  ( n8 ) & (n125 )  ;
assign n129 =  ( n128 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__97__ = n129 ;
assign __ILA_sha_acc_decode__[97] = __ILA_sha_decode_of_I__DOT__97__ ;
assign n130 =  ( n11 ) & (n125 )  ;
assign n131 =  ( n130 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__98__ = n131 ;
assign __ILA_sha_acc_decode__[98] = __ILA_sha_decode_of_I__DOT__98__ ;
assign n132 =  ( n14 ) & (n125 )  ;
assign n133 =  ( n132 ) & (n3 )  ;
assign __ILA_sha_decode_of_I__DOT__99__ = n133 ;
assign __ILA_sha_acc_decode__[99] = __ILA_sha_decode_of_I__DOT__99__ ;
assign n134 =  ( n126 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__100__ = n134 ;
assign __ILA_sha_acc_decode__[100] = __ILA_sha_decode_of_I__DOT__100__ ;
assign n135 =  ( n128 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__101__ = n135 ;
assign __ILA_sha_acc_decode__[101] = __ILA_sha_decode_of_I__DOT__101__ ;
assign n136 =  ( n130 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__102__ = n136 ;
assign __ILA_sha_acc_decode__[102] = __ILA_sha_decode_of_I__DOT__102__ ;
assign n137 =  ( n132 ) & (n17 )  ;
assign __ILA_sha_decode_of_I__DOT__103__ = n137 ;
assign __ILA_sha_acc_decode__[103] = __ILA_sha_decode_of_I__DOT__103__ ;
assign n138 =  ( n126 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__104__ = n138 ;
assign __ILA_sha_acc_decode__[104] = __ILA_sha_decode_of_I__DOT__104__ ;
assign n139 =  ( n128 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__105__ = n139 ;
assign __ILA_sha_acc_decode__[105] = __ILA_sha_decode_of_I__DOT__105__ ;
assign n140 =  ( n130 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__106__ = n140 ;
assign __ILA_sha_acc_decode__[106] = __ILA_sha_decode_of_I__DOT__106__ ;
assign n141 =  ( n132 ) & (n23 )  ;
assign __ILA_sha_decode_of_I__DOT__107__ = n141 ;
assign __ILA_sha_acc_decode__[107] = __ILA_sha_decode_of_I__DOT__107__ ;
assign n142 =  ( n126 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__108__ = n142 ;
assign __ILA_sha_acc_decode__[108] = __ILA_sha_decode_of_I__DOT__108__ ;
assign n143 =  ( n128 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__109__ = n143 ;
assign __ILA_sha_acc_decode__[109] = __ILA_sha_decode_of_I__DOT__109__ ;
assign n144 =  ( n130 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__110__ = n144 ;
assign __ILA_sha_acc_decode__[110] = __ILA_sha_decode_of_I__DOT__110__ ;
assign n145 =  ( n132 ) & (n29 )  ;
assign __ILA_sha_decode_of_I__DOT__111__ = n145 ;
assign __ILA_sha_acc_decode__[111] = __ILA_sha_decode_of_I__DOT__111__ ;
assign n146 =  ( n126 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__112__ = n146 ;
assign __ILA_sha_acc_decode__[112] = __ILA_sha_decode_of_I__DOT__112__ ;
assign n147 =  ( n128 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__113__ = n147 ;
assign __ILA_sha_acc_decode__[113] = __ILA_sha_decode_of_I__DOT__113__ ;
assign n148 =  ( n130 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__114__ = n148 ;
assign __ILA_sha_acc_decode__[114] = __ILA_sha_decode_of_I__DOT__114__ ;
assign n149 =  ( n132 ) & (n35 )  ;
assign __ILA_sha_decode_of_I__DOT__115__ = n149 ;
assign __ILA_sha_acc_decode__[115] = __ILA_sha_decode_of_I__DOT__115__ ;
assign n150 =  ( n126 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__116__ = n150 ;
assign __ILA_sha_acc_decode__[116] = __ILA_sha_decode_of_I__DOT__116__ ;
assign n151 =  ( n128 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__117__ = n151 ;
assign __ILA_sha_acc_decode__[117] = __ILA_sha_decode_of_I__DOT__117__ ;
assign n152 =  ( n130 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__118__ = n152 ;
assign __ILA_sha_acc_decode__[118] = __ILA_sha_decode_of_I__DOT__118__ ;
assign n153 =  ( n132 ) & (n41 )  ;
assign __ILA_sha_decode_of_I__DOT__119__ = n153 ;
assign __ILA_sha_acc_decode__[119] = __ILA_sha_decode_of_I__DOT__119__ ;
assign n154 =  ( n126 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__120__ = n154 ;
assign __ILA_sha_acc_decode__[120] = __ILA_sha_decode_of_I__DOT__120__ ;
assign n155 =  ( n128 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__121__ = n155 ;
assign __ILA_sha_acc_decode__[121] = __ILA_sha_decode_of_I__DOT__121__ ;
assign n156 =  ( n130 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__122__ = n156 ;
assign __ILA_sha_acc_decode__[122] = __ILA_sha_decode_of_I__DOT__122__ ;
assign n157 =  ( n132 ) & (n47 )  ;
assign __ILA_sha_decode_of_I__DOT__123__ = n157 ;
assign __ILA_sha_acc_decode__[123] = __ILA_sha_decode_of_I__DOT__123__ ;
assign n158 =  ( n126 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__124__ = n158 ;
assign __ILA_sha_acc_decode__[124] = __ILA_sha_decode_of_I__DOT__124__ ;
assign n159 =  ( n128 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__125__ = n159 ;
assign __ILA_sha_acc_decode__[125] = __ILA_sha_decode_of_I__DOT__125__ ;
assign n160 =  ( n130 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__126__ = n160 ;
assign __ILA_sha_acc_decode__[126] = __ILA_sha_decode_of_I__DOT__126__ ;
assign n161 =  ( n132 ) & (n53 )  ;
assign __ILA_sha_decode_of_I__DOT__127__ = n161 ;
assign __ILA_sha_acc_decode__[127] = __ILA_sha_decode_of_I__DOT__127__ ;
assign n162 =  ( n126 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__128__ = n162 ;
assign __ILA_sha_acc_decode__[128] = __ILA_sha_decode_of_I__DOT__128__ ;
assign n163 =  ( n128 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__129__ = n163 ;
assign __ILA_sha_acc_decode__[129] = __ILA_sha_decode_of_I__DOT__129__ ;
assign n164 =  ( n130 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__130__ = n164 ;
assign __ILA_sha_acc_decode__[130] = __ILA_sha_decode_of_I__DOT__130__ ;
assign n165 =  ( n132 ) & (n59 )  ;
assign __ILA_sha_decode_of_I__DOT__131__ = n165 ;
assign __ILA_sha_acc_decode__[131] = __ILA_sha_decode_of_I__DOT__131__ ;
assign n166 =  ( n126 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__132__ = n166 ;
assign __ILA_sha_acc_decode__[132] = __ILA_sha_decode_of_I__DOT__132__ ;
assign n167 =  ( n128 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__133__ = n167 ;
assign __ILA_sha_acc_decode__[133] = __ILA_sha_decode_of_I__DOT__133__ ;
assign n168 =  ( n130 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__134__ = n168 ;
assign __ILA_sha_acc_decode__[134] = __ILA_sha_decode_of_I__DOT__134__ ;
assign n169 =  ( n132 ) & (n65 )  ;
assign __ILA_sha_decode_of_I__DOT__135__ = n169 ;
assign __ILA_sha_acc_decode__[135] = __ILA_sha_decode_of_I__DOT__135__ ;
assign n170 =  ( n126 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__136__ = n170 ;
assign __ILA_sha_acc_decode__[136] = __ILA_sha_decode_of_I__DOT__136__ ;
assign n171 =  ( n128 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__137__ = n171 ;
assign __ILA_sha_acc_decode__[137] = __ILA_sha_decode_of_I__DOT__137__ ;
assign n172 =  ( n130 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__138__ = n172 ;
assign __ILA_sha_acc_decode__[138] = __ILA_sha_decode_of_I__DOT__138__ ;
assign n173 =  ( n132 ) & (n71 )  ;
assign __ILA_sha_decode_of_I__DOT__139__ = n173 ;
assign __ILA_sha_acc_decode__[139] = __ILA_sha_decode_of_I__DOT__139__ ;
assign n174 =  ( n126 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__140__ = n174 ;
assign __ILA_sha_acc_decode__[140] = __ILA_sha_decode_of_I__DOT__140__ ;
assign n175 =  ( n128 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__141__ = n175 ;
assign __ILA_sha_acc_decode__[141] = __ILA_sha_decode_of_I__DOT__141__ ;
assign n176 =  ( n130 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__142__ = n176 ;
assign __ILA_sha_acc_decode__[142] = __ILA_sha_decode_of_I__DOT__142__ ;
assign n177 =  ( n132 ) & (n77 )  ;
assign __ILA_sha_decode_of_I__DOT__143__ = n177 ;
assign __ILA_sha_acc_decode__[143] = __ILA_sha_decode_of_I__DOT__143__ ;
assign n178 =  ( n126 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__144__ = n178 ;
assign __ILA_sha_acc_decode__[144] = __ILA_sha_decode_of_I__DOT__144__ ;
assign n179 =  ( n128 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__145__ = n179 ;
assign __ILA_sha_acc_decode__[145] = __ILA_sha_decode_of_I__DOT__145__ ;
assign n180 =  ( n130 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__146__ = n180 ;
assign __ILA_sha_acc_decode__[146] = __ILA_sha_decode_of_I__DOT__146__ ;
assign n181 =  ( n132 ) & (n83 )  ;
assign __ILA_sha_decode_of_I__DOT__147__ = n181 ;
assign __ILA_sha_acc_decode__[147] = __ILA_sha_decode_of_I__DOT__147__ ;
assign n182 =  ( n126 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__148__ = n182 ;
assign __ILA_sha_acc_decode__[148] = __ILA_sha_decode_of_I__DOT__148__ ;
assign n183 =  ( n128 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__149__ = n183 ;
assign __ILA_sha_acc_decode__[149] = __ILA_sha_decode_of_I__DOT__149__ ;
assign n184 =  ( n130 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__150__ = n184 ;
assign __ILA_sha_acc_decode__[150] = __ILA_sha_decode_of_I__DOT__150__ ;
assign n185 =  ( n132 ) & (n89 )  ;
assign __ILA_sha_decode_of_I__DOT__151__ = n185 ;
assign __ILA_sha_acc_decode__[151] = __ILA_sha_decode_of_I__DOT__151__ ;
assign n186 =  ( n126 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__152__ = n186 ;
assign __ILA_sha_acc_decode__[152] = __ILA_sha_decode_of_I__DOT__152__ ;
assign n187 =  ( n128 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__153__ = n187 ;
assign __ILA_sha_acc_decode__[153] = __ILA_sha_decode_of_I__DOT__153__ ;
assign n188 =  ( n130 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__154__ = n188 ;
assign __ILA_sha_acc_decode__[154] = __ILA_sha_decode_of_I__DOT__154__ ;
assign n189 =  ( n132 ) & (n95 )  ;
assign __ILA_sha_decode_of_I__DOT__155__ = n189 ;
assign __ILA_sha_acc_decode__[155] = __ILA_sha_decode_of_I__DOT__155__ ;
assign n190 =  ( n126 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__156__ = n190 ;
assign __ILA_sha_acc_decode__[156] = __ILA_sha_decode_of_I__DOT__156__ ;
assign n191 =  ( n128 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__157__ = n191 ;
assign __ILA_sha_acc_decode__[157] = __ILA_sha_decode_of_I__DOT__157__ ;
assign n192 =  ( n130 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__158__ = n192 ;
assign __ILA_sha_acc_decode__[158] = __ILA_sha_decode_of_I__DOT__158__ ;
assign n193 =  ( n132 ) & (n101 )  ;
assign __ILA_sha_decode_of_I__DOT__159__ = n193 ;
assign __ILA_sha_acc_decode__[159] = __ILA_sha_decode_of_I__DOT__159__ ;
assign n194 =  ( sha_state ) == ( 3'd4 )  ;
assign n195 =  ( cmd ) == ( 2'd1 )  ;
assign n196 =  ( n194 ) & (n195 )  ;
assign n197 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n198 =  ( n196 ) & (n197 )  ;
assign n199 =  ( sha_state ) == ( 3'd3 )  ;
assign n200 =  ( cmd ) == ( 2'd1 )  ;
assign n201 =  ( n199 ) & (n200 )  ;
assign n202 =  ( n201 ) & (n197 )  ;
assign n203 =  ( sha_state ) == ( 3'd2 )  ;
assign n204 =  ( cmd ) == ( 2'd1 )  ;
assign n205 =  ( n203 ) & (n204 )  ;
assign n206 =  ( n205 ) & (n197 )  ;
assign n207 =  ( sha_state ) == ( 3'd1 )  ;
assign n208 =  ( cmd ) == ( 2'd1 )  ;
assign n209 =  ( n207 ) & (n208 )  ;
assign n210 =  ( n209 ) & (n197 )  ;
assign n211 =  ( sha_state ) == ( 3'd0 )  ;
assign n212 =  ( n211 ) & (n195 )  ;
assign n213 =  ( n212 ) & (n197 )  ;
assign n214 =  ( n210 ) | ( n213 )  ;
assign n215 =  ( n206 ) | ( n214 )  ;
assign n216 =  ( n202 ) | ( n215 )  ;
assign n217 =  ( n198 ) | ( n216 )  ;
assign n218 = sha_len[15:8] ;
assign n219 =  ( sha_state ) == ( 3'd4 )  ;
assign n220 =  ( cmd ) == ( 2'd1 )  ;
assign n221 =  ( n219 ) & (n220 )  ;
assign n222 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n223 =  ( n221 ) & (n222 )  ;
assign n224 =  ( sha_state ) == ( 3'd3 )  ;
assign n225 =  ( n224 ) & (n220 )  ;
assign n226 =  ( n225 ) & (n222 )  ;
assign n227 =  ( sha_state ) == ( 3'd2 )  ;
assign n228 =  ( n227 ) & (n220 )  ;
assign n229 =  ( n228 ) & (n222 )  ;
assign n230 =  ( sha_state ) == ( 3'd1 )  ;
assign n231 =  ( n230 ) & (n220 )  ;
assign n232 =  ( n231 ) & (n222 )  ;
assign n233 =  ( sha_state ) == ( 3'd0 )  ;
assign n234 =  ( n233 ) & (n220 )  ;
assign n235 =  ( n234 ) & (n222 )  ;
assign n236 =  ( n232 ) | ( n235 )  ;
assign n237 =  ( n229 ) | ( n236 )  ;
assign n238 =  ( n226 ) | ( n237 )  ;
assign n239 =  ( n223 ) | ( n238 )  ;
assign n240 = sha_len[7:0] ;
assign n241 =  ( sha_state ) == ( 3'd4 )  ;
assign n242 =  ( cmd ) == ( 2'd1 )  ;
assign n243 =  ( n241 ) & (n242 )  ;
assign n244 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n245 =  ( n243 ) & (n244 )  ;
assign n246 =  ( sha_state ) == ( 3'd3 )  ;
assign n247 =  ( n246 ) & (n242 )  ;
assign n248 =  ( n247 ) & (n244 )  ;
assign n249 =  ( sha_state ) == ( 3'd2 )  ;
assign n250 =  ( n249 ) & (n242 )  ;
assign n251 =  ( n250 ) & (n244 )  ;
assign n252 =  ( sha_state ) == ( 3'd1 )  ;
assign n253 =  ( n252 ) & (n242 )  ;
assign n254 =  ( n253 ) & (n244 )  ;
assign n255 =  ( sha_state ) == ( 3'd0 )  ;
assign n256 =  ( n255 ) & (n242 )  ;
assign n257 =  ( n256 ) & (n244 )  ;
assign n258 =  ( n254 ) | ( n257 )  ;
assign n259 =  ( n251 ) | ( n258 )  ;
assign n260 =  ( n248 ) | ( n259 )  ;
assign n261 =  ( n245 ) | ( n260 )  ;
assign n262 = sha_wraddr[15:8] ;
assign n263 =  ( sha_state ) == ( 3'd4 )  ;
assign n264 =  ( cmd ) == ( 2'd1 )  ;
assign n265 =  ( n263 ) & (n264 )  ;
assign n266 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n267 =  ( n265 ) & (n266 )  ;
assign n268 =  ( sha_state ) == ( 3'd3 )  ;
assign n269 =  ( n268 ) & (n264 )  ;
assign n270 =  ( n269 ) & (n266 )  ;
assign n271 =  ( sha_state ) == ( 3'd2 )  ;
assign n272 =  ( n271 ) & (n264 )  ;
assign n273 =  ( n272 ) & (n266 )  ;
assign n274 =  ( sha_state ) == ( 3'd1 )  ;
assign n275 =  ( n274 ) & (n264 )  ;
assign n276 =  ( n275 ) & (n266 )  ;
assign n277 =  ( sha_state ) == ( 3'd0 )  ;
assign n278 =  ( n277 ) & (n264 )  ;
assign n279 =  ( n278 ) & (n266 )  ;
assign n280 =  ( n276 ) | ( n279 )  ;
assign n281 =  ( n273 ) | ( n280 )  ;
assign n282 =  ( n270 ) | ( n281 )  ;
assign n283 =  ( n267 ) | ( n282 )  ;
assign n284 = sha_wraddr[7:0] ;
assign n285 =  ( sha_state ) == ( 3'd4 )  ;
assign n286 =  ( cmd ) == ( 2'd1 )  ;
assign n287 =  ( n285 ) & (n286 )  ;
assign n288 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n289 =  ( n287 ) & (n288 )  ;
assign n290 =  ( sha_state ) == ( 3'd3 )  ;
assign n291 =  ( n290 ) & (n286 )  ;
assign n292 =  ( n291 ) & (n288 )  ;
assign n293 =  ( sha_state ) == ( 3'd2 )  ;
assign n294 =  ( n293 ) & (n286 )  ;
assign n295 =  ( n294 ) & (n288 )  ;
assign n296 =  ( sha_state ) == ( 3'd1 )  ;
assign n297 =  ( n296 ) & (n286 )  ;
assign n298 =  ( n297 ) & (n288 )  ;
assign n299 =  ( sha_state ) == ( 3'd0 )  ;
assign n300 =  ( n299 ) & (n286 )  ;
assign n301 =  ( n300 ) & (n288 )  ;
assign n302 =  ( n298 ) | ( n301 )  ;
assign n303 =  ( n295 ) | ( n302 )  ;
assign n304 =  ( n292 ) | ( n303 )  ;
assign n305 =  ( n289 ) | ( n304 )  ;
assign n306 = sha_rdaddr[15:8] ;
assign n307 =  ( sha_state ) == ( 3'd4 )  ;
assign n308 =  ( cmd ) == ( 2'd1 )  ;
assign n309 =  ( n307 ) & (n308 )  ;
assign n310 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n311 =  ( n309 ) & (n310 )  ;
assign n312 =  ( sha_state ) == ( 3'd3 )  ;
assign n313 =  ( n312 ) & (n308 )  ;
assign n314 =  ( n313 ) & (n310 )  ;
assign n315 =  ( sha_state ) == ( 3'd2 )  ;
assign n316 =  ( n315 ) & (n308 )  ;
assign n317 =  ( n316 ) & (n310 )  ;
assign n318 =  ( sha_state ) == ( 3'd1 )  ;
assign n319 =  ( n318 ) & (n308 )  ;
assign n320 =  ( n319 ) & (n310 )  ;
assign n321 =  ( sha_state ) == ( 3'd0 )  ;
assign n322 =  ( n321 ) & (n308 )  ;
assign n323 =  ( n322 ) & (n310 )  ;
assign n324 =  ( n320 ) | ( n323 )  ;
assign n325 =  ( n317 ) | ( n324 )  ;
assign n326 =  ( n314 ) | ( n325 )  ;
assign n327 =  ( n311 ) | ( n326 )  ;
assign n328 = sha_rdaddr[7:0] ;
assign n329 =  ( cmd ) == ( 2'd2 )  ;
assign n330 =  ( n211 ) & (n329 )  ;
assign n331 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n332 =  ( n330 ) & (n331 )  ;
assign n333 =  ( sha_state ) == ( 3'd4 )  ;
assign n334 =  ( cmd ) == ( 2'd1 )  ;
assign n335 =  ( n333 ) & (n334 )  ;
assign n336 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n337 =  ( n335 ) & (n336 )  ;
assign n338 =  ( sha_state ) == ( 3'd3 )  ;
assign n339 =  ( n338 ) & (n334 )  ;
assign n340 =  ( n339 ) & (n336 )  ;
assign n341 =  ( sha_state ) == ( 3'd2 )  ;
assign n342 =  ( n341 ) & (n334 )  ;
assign n343 =  ( n342 ) & (n336 )  ;
assign n344 =  ( sha_state ) == ( 3'd1 )  ;
assign n345 =  ( n344 ) & (n334 )  ;
assign n346 =  ( n345 ) & (n336 )  ;
assign n347 =  ( n343 ) | ( n346 )  ;
assign n348 =  ( n340 ) | ( n347 )  ;
assign n349 =  ( n337 ) | ( n348 )  ;
assign n350 =  ( n332 ) | ( n349 )  ;
assign n351 =  {5'd0 , sha_state}  ;
assign n352 =  ( cmd ) == ( 2'd1 )  ;
assign n353 = ~ ( n352 )  ;
assign n354 =  ( n194 ) & (n353 )  ;
assign n355 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n356 =  ( n354 ) & (n355 )  ;
assign n357 =  ( cmd ) == ( 2'd1 )  ;
assign n358 = ~ ( n357 )  ;
assign n359 =  ( n199 ) & (n358 )  ;
assign n360 =  ( n359 ) & (n355 )  ;
assign n361 =  ( cmd ) == ( 2'd1 )  ;
assign n362 = ~ ( n361 )  ;
assign n363 =  ( n203 ) & (n362 )  ;
assign n364 =  ( n363 ) & (n355 )  ;
assign n365 = ~ ( n200 )  ;
assign n366 =  ( n207 ) & (n365 )  ;
assign n367 =  ( n366 ) & (n355 )  ;
assign n368 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n369 =  ( n354 ) & (n368 )  ;
assign n370 =  ( n359 ) & (n368 )  ;
assign n371 =  ( n363 ) & (n368 )  ;
assign n372 =  ( n366 ) & (n368 )  ;
assign n373 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n374 =  ( n354 ) & (n373 )  ;
assign n375 =  ( n359 ) & (n373 )  ;
assign n376 =  ( n363 ) & (n373 )  ;
assign n377 =  ( n366 ) & (n373 )  ;
assign n378 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n379 =  ( n354 ) & (n378 )  ;
assign n380 =  ( n359 ) & (n378 )  ;
assign n381 =  ( n363 ) & (n378 )  ;
assign n382 =  ( n366 ) & (n378 )  ;
assign n383 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n384 =  ( n354 ) & (n383 )  ;
assign n385 =  ( n359 ) & (n383 )  ;
assign n386 =  ( n363 ) & (n383 )  ;
assign n387 =  ( n366 ) & (n383 )  ;
assign n388 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n389 =  ( n354 ) & (n388 )  ;
assign n390 =  ( n359 ) & (n388 )  ;
assign n391 =  ( n363 ) & (n388 )  ;
assign n392 =  ( n366 ) & (n388 )  ;
assign n393 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n394 =  ( n354 ) & (n393 )  ;
assign n395 =  ( n359 ) & (n393 )  ;
assign n396 =  ( n363 ) & (n393 )  ;
assign n397 =  ( n366 ) & (n393 )  ;
assign n398 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n399 =  ( n354 ) & (n398 )  ;
assign n400 =  ( n359 ) & (n398 )  ;
assign n401 =  ( n363 ) & (n398 )  ;
assign n402 =  ( n366 ) & (n398 )  ;
assign n403 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n404 =  ( n354 ) & (n403 )  ;
assign n405 =  ( n359 ) & (n403 )  ;
assign n406 =  ( n363 ) & (n403 )  ;
assign n407 =  ( n366 ) & (n403 )  ;
assign n408 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n409 =  ( n354 ) & (n408 )  ;
assign n410 =  ( n359 ) & (n408 )  ;
assign n411 =  ( n363 ) & (n408 )  ;
assign n412 =  ( n366 ) & (n408 )  ;
assign n413 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n414 =  ( n354 ) & (n413 )  ;
assign n415 =  ( n359 ) & (n413 )  ;
assign n416 =  ( n363 ) & (n413 )  ;
assign n417 =  ( n366 ) & (n413 )  ;
assign n418 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n419 =  ( n354 ) & (n418 )  ;
assign n420 =  ( n359 ) & (n418 )  ;
assign n421 =  ( n363 ) & (n418 )  ;
assign n422 =  ( n366 ) & (n418 )  ;
assign n423 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n424 =  ( n354 ) & (n423 )  ;
assign n425 =  ( n359 ) & (n423 )  ;
assign n426 =  ( n363 ) & (n423 )  ;
assign n427 =  ( n366 ) & (n423 )  ;
assign n428 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n429 =  ( n354 ) & (n428 )  ;
assign n430 =  ( n359 ) & (n428 )  ;
assign n431 =  ( n363 ) & (n428 )  ;
assign n432 =  ( n366 ) & (n428 )  ;
assign n433 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n434 =  ( n354 ) & (n433 )  ;
assign n435 =  ( n359 ) & (n433 )  ;
assign n436 =  ( n363 ) & (n433 )  ;
assign n437 =  ( n366 ) & (n433 )  ;
assign n438 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n439 =  ( n354 ) & (n438 )  ;
assign n440 =  ( n359 ) & (n438 )  ;
assign n441 =  ( n363 ) & (n438 )  ;
assign n442 =  ( n366 ) & (n438 )  ;
assign n443 =  ( sha_state ) == ( 3'd0 )  ;
assign n444 =  ( cmd ) == ( 2'd2 )  ;
assign n445 =  ( n443 ) & (n444 )  ;
assign n446 =  ( n445 ) & (n355 )  ;
assign n447 =  ( n445 ) & (n368 )  ;
assign n448 =  ( n445 ) & (n373 )  ;
assign n449 =  ( n445 ) & (n378 )  ;
assign n450 =  ( n445 ) & (n383 )  ;
assign n451 =  ( n445 ) & (n388 )  ;
assign n452 =  ( n445 ) & (n393 )  ;
assign n453 =  ( n445 ) & (n398 )  ;
assign n454 =  ( n445 ) & (n403 )  ;
assign n455 =  ( n445 ) & (n408 )  ;
assign n456 =  ( n445 ) & (n413 )  ;
assign n457 =  ( n445 ) & (n418 )  ;
assign n458 =  ( n445 ) & (n428 )  ;
assign n459 =  ( n445 ) & (n433 )  ;
assign n460 =  ( n445 ) & (n438 )  ;
assign n461 =  ( sha_state ) == ( 3'd4 )  ;
assign n462 =  ( cmd ) == ( 2'd1 )  ;
assign n463 =  ( n461 ) & (n462 )  ;
assign n464 =  ( n463 ) & (n355 )  ;
assign n465 =  ( sha_state ) == ( 3'd3 )  ;
assign n466 =  ( n465 ) & (n462 )  ;
assign n467 =  ( n466 ) & (n355 )  ;
assign n468 =  ( sha_state ) == ( 3'd2 )  ;
assign n469 =  ( n468 ) & (n462 )  ;
assign n470 =  ( n469 ) & (n355 )  ;
assign n471 =  ( sha_state ) == ( 3'd1 )  ;
assign n472 =  ( n471 ) & (n462 )  ;
assign n473 =  ( n472 ) & (n355 )  ;
assign n474 =  ( sha_state ) == ( 3'd0 )  ;
assign n475 =  ( n474 ) & (n334 )  ;
assign n476 =  ( n475 ) & (n355 )  ;
assign n477 =  ( n463 ) & (n368 )  ;
assign n478 =  ( n466 ) & (n368 )  ;
assign n479 =  ( n469 ) & (n368 )  ;
assign n480 =  ( n472 ) & (n368 )  ;
assign n481 =  ( n475 ) & (n368 )  ;
assign n482 =  ( n463 ) & (n373 )  ;
assign n483 =  ( n466 ) & (n373 )  ;
assign n484 =  ( n469 ) & (n373 )  ;
assign n485 =  ( n472 ) & (n373 )  ;
assign n486 =  ( n475 ) & (n373 )  ;
assign n487 =  ( n463 ) & (n378 )  ;
assign n488 =  ( n466 ) & (n378 )  ;
assign n489 =  ( n469 ) & (n378 )  ;
assign n490 =  ( n472 ) & (n378 )  ;
assign n491 =  ( n475 ) & (n378 )  ;
assign n492 =  ( n463 ) & (n383 )  ;
assign n493 =  ( n466 ) & (n383 )  ;
assign n494 =  ( n469 ) & (n383 )  ;
assign n495 =  ( n472 ) & (n383 )  ;
assign n496 =  ( n475 ) & (n383 )  ;
assign n497 =  ( n463 ) & (n388 )  ;
assign n498 =  ( n466 ) & (n388 )  ;
assign n499 =  ( n469 ) & (n388 )  ;
assign n500 =  ( n472 ) & (n388 )  ;
assign n501 =  ( n475 ) & (n388 )  ;
assign n502 =  ( n463 ) & (n393 )  ;
assign n503 =  ( n466 ) & (n393 )  ;
assign n504 =  ( n469 ) & (n393 )  ;
assign n505 =  ( n472 ) & (n393 )  ;
assign n506 =  ( n475 ) & (n393 )  ;
assign n507 =  ( n463 ) & (n398 )  ;
assign n508 =  ( n466 ) & (n398 )  ;
assign n509 =  ( n469 ) & (n398 )  ;
assign n510 =  ( n472 ) & (n398 )  ;
assign n511 =  ( n475 ) & (n398 )  ;
assign n512 =  ( n475 ) & (n433 )  ;
assign n513 =  ( n463 ) & (n438 )  ;
assign n514 =  ( n466 ) & (n438 )  ;
assign n515 =  ( n469 ) & (n438 )  ;
assign n516 =  ( n472 ) & (n438 )  ;
assign n517 =  ( n475 ) & (n438 )  ;
assign n518 =  ( n516 ) | ( n517 )  ;
assign n519 =  ( n515 ) | ( n518 )  ;
assign n520 =  ( n514 ) | ( n519 )  ;
assign n521 =  ( n513 ) | ( n520 )  ;
assign n522 =  ( n512 ) | ( n521 )  ;
assign n523 =  ( n511 ) | ( n522 )  ;
assign n524 =  ( n510 ) | ( n523 )  ;
assign n525 =  ( n509 ) | ( n524 )  ;
assign n526 =  ( n508 ) | ( n525 )  ;
assign n527 =  ( n507 ) | ( n526 )  ;
assign n528 =  ( n506 ) | ( n527 )  ;
assign n529 =  ( n505 ) | ( n528 )  ;
assign n530 =  ( n504 ) | ( n529 )  ;
assign n531 =  ( n503 ) | ( n530 )  ;
assign n532 =  ( n502 ) | ( n531 )  ;
assign n533 =  ( n501 ) | ( n532 )  ;
assign n534 =  ( n500 ) | ( n533 )  ;
assign n535 =  ( n499 ) | ( n534 )  ;
assign n536 =  ( n498 ) | ( n535 )  ;
assign n537 =  ( n497 ) | ( n536 )  ;
assign n538 =  ( n496 ) | ( n537 )  ;
assign n539 =  ( n495 ) | ( n538 )  ;
assign n540 =  ( n494 ) | ( n539 )  ;
assign n541 =  ( n493 ) | ( n540 )  ;
assign n542 =  ( n492 ) | ( n541 )  ;
assign n543 =  ( n491 ) | ( n542 )  ;
assign n544 =  ( n490 ) | ( n543 )  ;
assign n545 =  ( n489 ) | ( n544 )  ;
assign n546 =  ( n488 ) | ( n545 )  ;
assign n547 =  ( n487 ) | ( n546 )  ;
assign n548 =  ( n486 ) | ( n547 )  ;
assign n549 =  ( n485 ) | ( n548 )  ;
assign n550 =  ( n484 ) | ( n549 )  ;
assign n551 =  ( n483 ) | ( n550 )  ;
assign n552 =  ( n482 ) | ( n551 )  ;
assign n553 =  ( n481 ) | ( n552 )  ;
assign n554 =  ( n480 ) | ( n553 )  ;
assign n555 =  ( n479 ) | ( n554 )  ;
assign n556 =  ( n478 ) | ( n555 )  ;
assign n557 =  ( n477 ) | ( n556 )  ;
assign n558 =  ( n476 ) | ( n557 )  ;
assign n559 =  ( n473 ) | ( n558 )  ;
assign n560 =  ( n470 ) | ( n559 )  ;
assign n561 =  ( n467 ) | ( n560 )  ;
assign n562 =  ( n464 ) | ( n561 )  ;
assign n563 =  ( n460 ) | ( n562 )  ;
assign n564 =  ( n459 ) | ( n563 )  ;
assign n565 =  ( n458 ) | ( n564 )  ;
assign n566 =  ( n457 ) | ( n565 )  ;
assign n567 =  ( n456 ) | ( n566 )  ;
assign n568 =  ( n455 ) | ( n567 )  ;
assign n569 =  ( n454 ) | ( n568 )  ;
assign n570 =  ( n453 ) | ( n569 )  ;
assign n571 =  ( n452 ) | ( n570 )  ;
assign n572 =  ( n451 ) | ( n571 )  ;
assign n573 =  ( n450 ) | ( n572 )  ;
assign n574 =  ( n449 ) | ( n573 )  ;
assign n575 =  ( n448 ) | ( n574 )  ;
assign n576 =  ( n447 ) | ( n575 )  ;
assign n577 =  ( n446 ) | ( n576 )  ;
assign n578 =  ( n442 ) | ( n577 )  ;
assign n579 =  ( n441 ) | ( n578 )  ;
assign n580 =  ( n440 ) | ( n579 )  ;
assign n581 =  ( n439 ) | ( n580 )  ;
assign n582 =  ( n437 ) | ( n581 )  ;
assign n583 =  ( n436 ) | ( n582 )  ;
assign n584 =  ( n435 ) | ( n583 )  ;
assign n585 =  ( n434 ) | ( n584 )  ;
assign n586 =  ( n432 ) | ( n585 )  ;
assign n587 =  ( n431 ) | ( n586 )  ;
assign n588 =  ( n430 ) | ( n587 )  ;
assign n589 =  ( n429 ) | ( n588 )  ;
assign n590 =  ( n427 ) | ( n589 )  ;
assign n591 =  ( n426 ) | ( n590 )  ;
assign n592 =  ( n425 ) | ( n591 )  ;
assign n593 =  ( n424 ) | ( n592 )  ;
assign n594 =  ( n422 ) | ( n593 )  ;
assign n595 =  ( n421 ) | ( n594 )  ;
assign n596 =  ( n420 ) | ( n595 )  ;
assign n597 =  ( n419 ) | ( n596 )  ;
assign n598 =  ( n417 ) | ( n597 )  ;
assign n599 =  ( n416 ) | ( n598 )  ;
assign n600 =  ( n415 ) | ( n599 )  ;
assign n601 =  ( n414 ) | ( n600 )  ;
assign n602 =  ( n412 ) | ( n601 )  ;
assign n603 =  ( n411 ) | ( n602 )  ;
assign n604 =  ( n410 ) | ( n603 )  ;
assign n605 =  ( n409 ) | ( n604 )  ;
assign n606 =  ( n407 ) | ( n605 )  ;
assign n607 =  ( n406 ) | ( n606 )  ;
assign n608 =  ( n405 ) | ( n607 )  ;
assign n609 =  ( n404 ) | ( n608 )  ;
assign n610 =  ( n402 ) | ( n609 )  ;
assign n611 =  ( n401 ) | ( n610 )  ;
assign n612 =  ( n400 ) | ( n611 )  ;
assign n613 =  ( n399 ) | ( n612 )  ;
assign n614 =  ( n397 ) | ( n613 )  ;
assign n615 =  ( n396 ) | ( n614 )  ;
assign n616 =  ( n395 ) | ( n615 )  ;
assign n617 =  ( n394 ) | ( n616 )  ;
assign n618 =  ( n392 ) | ( n617 )  ;
assign n619 =  ( n391 ) | ( n618 )  ;
assign n620 =  ( n390 ) | ( n619 )  ;
assign n621 =  ( n389 ) | ( n620 )  ;
assign n622 =  ( n387 ) | ( n621 )  ;
assign n623 =  ( n386 ) | ( n622 )  ;
assign n624 =  ( n385 ) | ( n623 )  ;
assign n625 =  ( n384 ) | ( n624 )  ;
assign n626 =  ( n382 ) | ( n625 )  ;
assign n627 =  ( n381 ) | ( n626 )  ;
assign n628 =  ( n380 ) | ( n627 )  ;
assign n629 =  ( n379 ) | ( n628 )  ;
assign n630 =  ( n377 ) | ( n629 )  ;
assign n631 =  ( n376 ) | ( n630 )  ;
assign n632 =  ( n375 ) | ( n631 )  ;
assign n633 =  ( n374 ) | ( n632 )  ;
assign n634 =  ( n372 ) | ( n633 )  ;
assign n635 =  ( n371 ) | ( n634 )  ;
assign n636 =  ( n370 ) | ( n635 )  ;
assign n637 =  ( n369 ) | ( n636 )  ;
assign n638 =  ( n367 ) | ( n637 )  ;
assign n639 =  ( n364 ) | ( n638 )  ;
assign n640 =  ( n360 ) | ( n639 )  ;
assign n641 =  ( n356 ) | ( n640 )  ;
assign n642 =  ( n641 ) ? ( 8'd0 ) : ( dataout ) ;
assign n643 =  ( n350 ) ? ( n351 ) : ( n642 ) ;
assign n644 =  ( n327 ) ? ( n328 ) : ( n643 ) ;
assign n645 =  ( n305 ) ? ( n306 ) : ( n644 ) ;
assign n646 =  ( n283 ) ? ( n284 ) : ( n645 ) ;
assign n647 =  ( n261 ) ? ( n262 ) : ( n646 ) ;
assign n648 =  ( n239 ) ? ( n240 ) : ( n647 ) ;
assign n649 =  ( n217 ) ? ( n218 ) : ( n648 ) ;
assign n650 =  ( sha_state ) == ( 3'd1 )  ;
assign n651 = ~ ( n195 )  ;
assign n652 =  ( n650 ) & (n651 )  ;
assign n653 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n654 =  ( n652 ) & (n653 )  ;
assign n655 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n656 =  ( n652 ) & (n655 )  ;
assign n657 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n658 =  ( n652 ) & (n657 )  ;
assign n659 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n660 =  ( n652 ) & (n659 )  ;
assign n661 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n662 =  ( n652 ) & (n661 )  ;
assign n663 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n664 =  ( n652 ) & (n663 )  ;
assign n665 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n666 =  ( n652 ) & (n665 )  ;
assign n667 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n668 =  ( n652 ) & (n667 )  ;
assign n669 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n670 =  ( n652 ) & (n669 )  ;
assign n671 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n672 =  ( n652 ) & (n671 )  ;
assign n673 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n674 =  ( n652 ) & (n673 )  ;
assign n675 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n676 =  ( n652 ) & (n675 )  ;
assign n677 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n678 =  ( n652 ) & (n677 )  ;
assign n679 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n680 =  ( n652 ) & (n679 )  ;
assign n681 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n682 =  ( n652 ) & (n681 )  ;
assign n683 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n684 =  ( n652 ) & (n683 )  ;
assign n685 =  ( n650 ) & (n357 )  ;
assign n686 =  ( n685 ) & (n653 )  ;
assign n687 =  ( n685 ) & (n655 )  ;
assign n688 =  ( n685 ) & (n657 )  ;
assign n689 =  ( n685 ) & (n659 )  ;
assign n690 =  ( n685 ) & (n661 )  ;
assign n691 =  ( n685 ) & (n663 )  ;
assign n692 =  ( n685 ) & (n665 )  ;
assign n693 =  ( n685 ) & (n667 )  ;
assign n694 =  ( n685 ) & (n669 )  ;
assign n695 =  ( n685 ) & (n671 )  ;
assign n696 =  ( n685 ) & (n673 )  ;
assign n697 =  ( n685 ) & (n675 )  ;
assign n698 =  ( n685 ) & (n677 )  ;
assign n699 =  ( n685 ) & (n679 )  ;
assign n700 =  ( n685 ) & (n681 )  ;
assign n701 =  ( n685 ) & (n683 )  ;
assign n702 =  ( n700 ) | ( n701 )  ;
assign n703 =  ( n699 ) | ( n702 )  ;
assign n704 =  ( n698 ) | ( n703 )  ;
assign n705 =  ( n697 ) | ( n704 )  ;
assign n706 =  ( n696 ) | ( n705 )  ;
assign n707 =  ( n695 ) | ( n706 )  ;
assign n708 =  ( n694 ) | ( n707 )  ;
assign n709 =  ( n693 ) | ( n708 )  ;
assign n710 =  ( n692 ) | ( n709 )  ;
assign n711 =  ( n691 ) | ( n710 )  ;
assign n712 =  ( n690 ) | ( n711 )  ;
assign n713 =  ( n689 ) | ( n712 )  ;
assign n714 =  ( n688 ) | ( n713 )  ;
assign n715 =  ( n687 ) | ( n714 )  ;
assign n716 =  ( n686 ) | ( n715 )  ;
assign n717 =  ( n684 ) | ( n716 )  ;
assign n718 =  ( n682 ) | ( n717 )  ;
assign n719 =  ( n680 ) | ( n718 )  ;
assign n720 =  ( n678 ) | ( n719 )  ;
assign n721 =  ( n676 ) | ( n720 )  ;
assign n722 =  ( n674 ) | ( n721 )  ;
assign n723 =  ( n672 ) | ( n722 )  ;
assign n724 =  ( n670 ) | ( n723 )  ;
assign n725 =  ( n668 ) | ( n724 )  ;
assign n726 =  ( n666 ) | ( n725 )  ;
assign n727 =  ( n664 ) | ( n726 )  ;
assign n728 =  ( n662 ) | ( n727 )  ;
assign n729 =  ( n660 ) | ( n728 )  ;
assign n730 =  ( n658 ) | ( n729 )  ;
assign n731 =  ( n656 ) | ( n730 )  ;
assign n732 =  ( n654 ) | ( n731 )  ;
assign n733 =  ( sha_bytes_read ) + ( 16'd64 )  ;
assign n734 =  ( n732 ) ? ( n733 ) : ( sha_bytes_read ) ;
assign n735 =  ( cmddata ) == ( 8'd1 )  ;
assign n736 =  ( n735 ) ? ( 16'd0 ) : ( sha_bytes_read ) ;
assign n737 =  ( sha_state ) == ( 3'd3 )  ;
assign n738 =  ( cmd ) == ( 2'd1 )  ;
assign n739 = ~ ( n738 )  ;
assign n740 =  ( n737 ) & (n739 )  ;
assign n741 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n742 =  ( n740 ) & (n741 )  ;
assign n743 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n744 =  ( n740 ) & (n743 )  ;
assign n745 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n746 =  ( n740 ) & (n745 )  ;
assign n747 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n748 =  ( n740 ) & (n747 )  ;
assign n749 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n750 =  ( n740 ) & (n749 )  ;
assign n751 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n752 =  ( n740 ) & (n751 )  ;
assign n753 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n754 =  ( n740 ) & (n753 )  ;
assign n755 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n756 =  ( n740 ) & (n755 )  ;
assign n757 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n758 =  ( n740 ) & (n757 )  ;
assign n759 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n760 =  ( n740 ) & (n759 )  ;
assign n761 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n762 =  ( n740 ) & (n761 )  ;
assign n763 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n764 =  ( n740 ) & (n763 )  ;
assign n765 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n766 =  ( n740 ) & (n765 )  ;
assign n767 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n768 =  ( n740 ) & (n767 )  ;
assign n769 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n770 =  ( n740 ) & (n769 )  ;
assign n771 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n772 =  ( n740 ) & (n771 )  ;
assign n773 =  ( n737 ) & (n361 )  ;
assign n774 =  ( n773 ) & (n741 )  ;
assign n775 =  ( n773 ) & (n743 )  ;
assign n776 =  ( n773 ) & (n745 )  ;
assign n777 =  ( n773 ) & (n747 )  ;
assign n778 =  ( n773 ) & (n749 )  ;
assign n779 =  ( n773 ) & (n751 )  ;
assign n780 =  ( n773 ) & (n753 )  ;
assign n781 =  ( n773 ) & (n755 )  ;
assign n782 =  ( n773 ) & (n757 )  ;
assign n783 =  ( n773 ) & (n759 )  ;
assign n784 =  ( n773 ) & (n761 )  ;
assign n785 =  ( n773 ) & (n763 )  ;
assign n786 =  ( n773 ) & (n765 )  ;
assign n787 =  ( n773 ) & (n767 )  ;
assign n788 =  ( n773 ) & (n769 )  ;
assign n789 =  ( n773 ) & (n771 )  ;
assign n790 =  ( n788 ) | ( n789 )  ;
assign n791 =  ( n787 ) | ( n790 )  ;
assign n792 =  ( n786 ) | ( n791 )  ;
assign n793 =  ( n785 ) | ( n792 )  ;
assign n794 =  ( n784 ) | ( n793 )  ;
assign n795 =  ( n783 ) | ( n794 )  ;
assign n796 =  ( n782 ) | ( n795 )  ;
assign n797 =  ( n781 ) | ( n796 )  ;
assign n798 =  ( n780 ) | ( n797 )  ;
assign n799 =  ( n779 ) | ( n798 )  ;
assign n800 =  ( n778 ) | ( n799 )  ;
assign n801 =  ( n777 ) | ( n800 )  ;
assign n802 =  ( n776 ) | ( n801 )  ;
assign n803 =  ( n775 ) | ( n802 )  ;
assign n804 =  ( n774 ) | ( n803 )  ;
assign n805 =  ( n772 ) | ( n804 )  ;
assign n806 =  ( n770 ) | ( n805 )  ;
assign n807 =  ( n768 ) | ( n806 )  ;
assign n808 =  ( n766 ) | ( n807 )  ;
assign n809 =  ( n764 ) | ( n808 )  ;
assign n810 =  ( n762 ) | ( n809 )  ;
assign n811 =  ( n760 ) | ( n810 )  ;
assign n812 =  ( n758 ) | ( n811 )  ;
assign n813 =  ( n756 ) | ( n812 )  ;
assign n814 =  ( n754 ) | ( n813 )  ;
assign n815 =  ( n752 ) | ( n814 )  ;
assign n816 =  ( n750 ) | ( n815 )  ;
assign n817 =  ( n748 ) | ( n816 )  ;
assign n818 =  ( n746 ) | ( n817 )  ;
assign n819 =  ( n744 ) | ( n818 )  ;
assign n820 =  ( n742 ) | ( n819 )  ;
fun_sha  applyFunc_n822(
    .arg0( sha_rd_data ),
    .result( n821 )
);
assign n823 = n821 ;
assign n824 =  ( n820 ) ? ( n823 ) : ( sha_hs_data ) ;
assign n825 = sha_len[15:8] ;
assign n826 =  { ( n825 ) , ( cmddata ) }  ;
assign n827 = sha_len[7:0] ;
assign n828 =  { ( cmddata ) , ( n827 ) }  ;
assign n829 =  ( sha_state ) == ( 3'd1 )  ;
assign n830 = ~ ( n204 )  ;
assign n831 =  ( n829 ) & (n830 )  ;
assign n832 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n833 =  ( n831 ) & (n832 )  ;
assign n834 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n835 =  ( n831 ) & (n834 )  ;
assign n836 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n837 =  ( n831 ) & (n836 )  ;
assign n838 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n839 =  ( n831 ) & (n838 )  ;
assign n840 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n841 =  ( n831 ) & (n840 )  ;
assign n842 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n843 =  ( n831 ) & (n842 )  ;
assign n844 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n845 =  ( n831 ) & (n844 )  ;
assign n846 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n847 =  ( n831 ) & (n846 )  ;
assign n848 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n849 =  ( n831 ) & (n848 )  ;
assign n850 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n851 =  ( n831 ) & (n850 )  ;
assign n852 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n853 =  ( n831 ) & (n852 )  ;
assign n854 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n855 =  ( n831 ) & (n854 )  ;
assign n856 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n857 =  ( n831 ) & (n856 )  ;
assign n858 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n859 =  ( n831 ) & (n858 )  ;
assign n860 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n861 =  ( n831 ) & (n860 )  ;
assign n862 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n863 =  ( n831 ) & (n862 )  ;
assign n864 =  ( n829 ) & (n352 )  ;
assign n865 =  ( n864 ) & (n832 )  ;
assign n866 =  ( n864 ) & (n834 )  ;
assign n867 =  ( n864 ) & (n836 )  ;
assign n868 =  ( n864 ) & (n838 )  ;
assign n869 =  ( n864 ) & (n840 )  ;
assign n870 =  ( n864 ) & (n842 )  ;
assign n871 =  ( n864 ) & (n844 )  ;
assign n872 =  ( n864 ) & (n846 )  ;
assign n873 =  ( n864 ) & (n848 )  ;
assign n874 =  ( n864 ) & (n850 )  ;
assign n875 =  ( n864 ) & (n852 )  ;
assign n876 =  ( n864 ) & (n854 )  ;
assign n877 =  ( n864 ) & (n856 )  ;
assign n878 =  ( n864 ) & (n858 )  ;
assign n879 =  ( n864 ) & (n860 )  ;
assign n880 =  ( n864 ) & (n862 )  ;
assign n881 =  ( n879 ) | ( n880 )  ;
assign n882 =  ( n878 ) | ( n881 )  ;
assign n883 =  ( n877 ) | ( n882 )  ;
assign n884 =  ( n876 ) | ( n883 )  ;
assign n885 =  ( n875 ) | ( n884 )  ;
assign n886 =  ( n874 ) | ( n885 )  ;
assign n887 =  ( n873 ) | ( n886 )  ;
assign n888 =  ( n872 ) | ( n887 )  ;
assign n889 =  ( n871 ) | ( n888 )  ;
assign n890 =  ( n870 ) | ( n889 )  ;
assign n891 =  ( n869 ) | ( n890 )  ;
assign n892 =  ( n868 ) | ( n891 )  ;
assign n893 =  ( n867 ) | ( n892 )  ;
assign n894 =  ( n866 ) | ( n893 )  ;
assign n895 =  ( n865 ) | ( n894 )  ;
assign n896 =  ( n863 ) | ( n895 )  ;
assign n897 =  ( n861 ) | ( n896 )  ;
assign n898 =  ( n859 ) | ( n897 )  ;
assign n899 =  ( n857 ) | ( n898 )  ;
assign n900 =  ( n855 ) | ( n899 )  ;
assign n901 =  ( n853 ) | ( n900 )  ;
assign n902 =  ( n851 ) | ( n901 )  ;
assign n903 =  ( n849 ) | ( n902 )  ;
assign n904 =  ( n847 ) | ( n903 )  ;
assign n905 =  ( n845 ) | ( n904 )  ;
assign n906 =  ( n843 ) | ( n905 )  ;
assign n907 =  ( n841 ) | ( n906 )  ;
assign n908 =  ( n839 ) | ( n907 )  ;
assign n909 =  ( n837 ) | ( n908 )  ;
assign n910 =  ( n835 ) | ( n909 )  ;
assign n911 =  ( n833 ) | ( n910 )  ;
assign n912 =  ( sha_rdaddr ) + ( sha_bytes_read )  ;
assign n913 =  ( n912 ) + ( 16'd0 )  ;
assign XRAM_addr_n914 = n913 ;
assign n916 = XRAM_data_n915 ;
assign n917 =  ( n912 ) + ( 16'd1 )  ;
assign XRAM_addr_n918 = n917 ;
assign n920 = XRAM_data_n919 ;
assign n921 =  { ( n916 ) , ( n920 ) }  ;
assign n922 =  ( n912 ) + ( 16'd2 )  ;
assign XRAM_addr_n923 = n922 ;
assign n925 = XRAM_data_n924 ;
assign n926 =  { ( n921 ) , ( n925 ) }  ;
assign n927 =  ( n912 ) + ( 16'd3 )  ;
assign XRAM_addr_n928 = n927 ;
assign n930 = XRAM_data_n929 ;
assign n931 =  { ( n926 ) , ( n930 ) }  ;
assign n932 =  ( n912 ) + ( 16'd4 )  ;
assign XRAM_addr_n933 = n932 ;
assign n935 = XRAM_data_n934 ;
assign n936 =  { ( n931 ) , ( n935 ) }  ;
assign n937 =  ( n912 ) + ( 16'd5 )  ;
assign XRAM_addr_n938 = n937 ;
assign n940 = XRAM_data_n939 ;
assign n941 =  { ( n936 ) , ( n940 ) }  ;
assign n942 =  ( n912 ) + ( 16'd6 )  ;
assign XRAM_addr_n943 = n942 ;
assign n945 = XRAM_data_n944 ;
assign n946 =  { ( n941 ) , ( n945 ) }  ;
assign n947 =  ( n912 ) + ( 16'd7 )  ;
assign XRAM_addr_n948 = n947 ;
assign n950 = XRAM_data_n949 ;
assign n951 =  { ( n946 ) , ( n950 ) }  ;
assign n952 =  ( n912 ) + ( 16'd8 )  ;
assign XRAM_addr_n953 = n952 ;
assign n955 = XRAM_data_n954 ;
assign n956 =  { ( n951 ) , ( n955 ) }  ;
assign n957 =  ( n912 ) + ( 16'd9 )  ;
assign XRAM_addr_n958 = n957 ;
assign n960 = XRAM_data_n959 ;
assign n961 =  { ( n956 ) , ( n960 ) }  ;
assign n962 =  ( n912 ) + ( 16'd10 )  ;
assign XRAM_addr_n963 = n962 ;
assign n965 = XRAM_data_n964 ;
assign n966 =  { ( n961 ) , ( n965 ) }  ;
assign n967 =  ( n912 ) + ( 16'd11 )  ;
assign XRAM_addr_n968 = n967 ;
assign n970 = XRAM_data_n969 ;
assign n971 =  { ( n966 ) , ( n970 ) }  ;
assign n972 =  ( n912 ) + ( 16'd12 )  ;
assign XRAM_addr_n973 = n972 ;
assign n975 = XRAM_data_n974 ;
assign n976 =  { ( n971 ) , ( n975 ) }  ;
assign n977 =  ( n912 ) + ( 16'd13 )  ;
assign XRAM_addr_n978 = n977 ;
assign n980 = XRAM_data_n979 ;
assign n981 =  { ( n976 ) , ( n980 ) }  ;
assign n982 =  ( n912 ) + ( 16'd14 )  ;
assign XRAM_addr_n983 = n982 ;
assign n985 = XRAM_data_n984 ;
assign n986 =  { ( n981 ) , ( n985 ) }  ;
assign n987 =  ( n912 ) + ( 16'd15 )  ;
assign XRAM_addr_n988 = n987 ;
assign n990 = XRAM_data_n989 ;
assign n991 =  { ( n986 ) , ( n990 ) }  ;
assign n992 =  ( n912 ) + ( 16'd16 )  ;
assign XRAM_addr_n993 = n992 ;
assign n995 = XRAM_data_n994 ;
assign n996 =  { ( n991 ) , ( n995 ) }  ;
assign n997 =  ( n912 ) + ( 16'd17 )  ;
assign XRAM_addr_n998 = n997 ;
assign n1000 = XRAM_data_n999 ;
assign n1001 =  { ( n996 ) , ( n1000 ) }  ;
assign n1002 =  ( n912 ) + ( 16'd18 )  ;
assign XRAM_addr_n1003 = n1002 ;
assign n1005 = XRAM_data_n1004 ;
assign n1006 =  { ( n1001 ) , ( n1005 ) }  ;
assign n1007 =  ( n912 ) + ( 16'd19 )  ;
assign XRAM_addr_n1008 = n1007 ;
assign n1010 = XRAM_data_n1009 ;
assign n1011 =  { ( n1006 ) , ( n1010 ) }  ;
assign n1012 =  ( n912 ) + ( 16'd20 )  ;
assign XRAM_addr_n1013 = n1012 ;
assign n1015 = XRAM_data_n1014 ;
assign n1016 =  { ( n1011 ) , ( n1015 ) }  ;
assign n1017 =  ( n912 ) + ( 16'd21 )  ;
assign XRAM_addr_n1018 = n1017 ;
assign n1020 = XRAM_data_n1019 ;
assign n1021 =  { ( n1016 ) , ( n1020 ) }  ;
assign n1022 =  ( n912 ) + ( 16'd22 )  ;
assign XRAM_addr_n1023 = n1022 ;
assign n1025 = XRAM_data_n1024 ;
assign n1026 =  { ( n1021 ) , ( n1025 ) }  ;
assign n1027 =  ( n912 ) + ( 16'd23 )  ;
assign XRAM_addr_n1028 = n1027 ;
assign n1030 = XRAM_data_n1029 ;
assign n1031 =  { ( n1026 ) , ( n1030 ) }  ;
assign n1032 =  ( n912 ) + ( 16'd24 )  ;
assign XRAM_addr_n1033 = n1032 ;
assign n1035 = XRAM_data_n1034 ;
assign n1036 =  { ( n1031 ) , ( n1035 ) }  ;
assign n1037 =  ( n912 ) + ( 16'd25 )  ;
assign XRAM_addr_n1038 = n1037 ;
assign n1040 = XRAM_data_n1039 ;
assign n1041 =  { ( n1036 ) , ( n1040 ) }  ;
assign n1042 =  ( n912 ) + ( 16'd26 )  ;
assign XRAM_addr_n1043 = n1042 ;
assign n1045 = XRAM_data_n1044 ;
assign n1046 =  { ( n1041 ) , ( n1045 ) }  ;
assign n1047 =  ( n912 ) + ( 16'd27 )  ;
assign XRAM_addr_n1048 = n1047 ;
assign n1050 = XRAM_data_n1049 ;
assign n1051 =  { ( n1046 ) , ( n1050 ) }  ;
assign n1052 =  ( n912 ) + ( 16'd28 )  ;
assign XRAM_addr_n1053 = n1052 ;
assign n1055 = XRAM_data_n1054 ;
assign n1056 =  { ( n1051 ) , ( n1055 ) }  ;
assign n1057 =  ( n912 ) + ( 16'd29 )  ;
assign XRAM_addr_n1058 = n1057 ;
assign n1060 = XRAM_data_n1059 ;
assign n1061 =  { ( n1056 ) , ( n1060 ) }  ;
assign n1062 =  ( n912 ) + ( 16'd30 )  ;
assign XRAM_addr_n1063 = n1062 ;
assign n1065 = XRAM_data_n1064 ;
assign n1066 =  { ( n1061 ) , ( n1065 ) }  ;
assign n1067 =  ( n912 ) + ( 16'd31 )  ;
assign XRAM_addr_n1068 = n1067 ;
assign n1070 = XRAM_data_n1069 ;
assign n1071 =  { ( n1066 ) , ( n1070 ) }  ;
assign n1072 =  ( n912 ) + ( 16'd32 )  ;
assign XRAM_addr_n1073 = n1072 ;
assign n1075 = XRAM_data_n1074 ;
assign n1076 =  { ( n1071 ) , ( n1075 ) }  ;
assign n1077 =  ( n912 ) + ( 16'd33 )  ;
assign XRAM_addr_n1078 = n1077 ;
assign n1080 = XRAM_data_n1079 ;
assign n1081 =  { ( n1076 ) , ( n1080 ) }  ;
assign n1082 =  ( n912 ) + ( 16'd34 )  ;
assign XRAM_addr_n1083 = n1082 ;
assign n1085 = XRAM_data_n1084 ;
assign n1086 =  { ( n1081 ) , ( n1085 ) }  ;
assign n1087 =  ( n912 ) + ( 16'd35 )  ;
assign XRAM_addr_n1088 = n1087 ;
assign n1090 = XRAM_data_n1089 ;
assign n1091 =  { ( n1086 ) , ( n1090 ) }  ;
assign n1092 =  ( n912 ) + ( 16'd36 )  ;
assign XRAM_addr_n1093 = n1092 ;
assign n1095 = XRAM_data_n1094 ;
assign n1096 =  { ( n1091 ) , ( n1095 ) }  ;
assign n1097 =  ( n912 ) + ( 16'd37 )  ;
assign XRAM_addr_n1098 = n1097 ;
assign n1100 = XRAM_data_n1099 ;
assign n1101 =  { ( n1096 ) , ( n1100 ) }  ;
assign n1102 =  ( n912 ) + ( 16'd38 )  ;
assign XRAM_addr_n1103 = n1102 ;
assign n1105 = XRAM_data_n1104 ;
assign n1106 =  { ( n1101 ) , ( n1105 ) }  ;
assign n1107 =  ( n912 ) + ( 16'd39 )  ;
assign XRAM_addr_n1108 = n1107 ;
assign n1110 = XRAM_data_n1109 ;
assign n1111 =  { ( n1106 ) , ( n1110 ) }  ;
assign n1112 =  ( n912 ) + ( 16'd40 )  ;
assign XRAM_addr_n1113 = n1112 ;
assign n1115 = XRAM_data_n1114 ;
assign n1116 =  { ( n1111 ) , ( n1115 ) }  ;
assign n1117 =  ( n912 ) + ( 16'd41 )  ;
assign XRAM_addr_n1118 = n1117 ;
assign n1120 = XRAM_data_n1119 ;
assign n1121 =  { ( n1116 ) , ( n1120 ) }  ;
assign n1122 =  ( n912 ) + ( 16'd42 )  ;
assign XRAM_addr_n1123 = n1122 ;
assign n1125 = XRAM_data_n1124 ;
assign n1126 =  { ( n1121 ) , ( n1125 ) }  ;
assign n1127 =  ( n912 ) + ( 16'd43 )  ;
assign XRAM_addr_n1128 = n1127 ;
assign n1130 = XRAM_data_n1129 ;
assign n1131 =  { ( n1126 ) , ( n1130 ) }  ;
assign n1132 =  ( n912 ) + ( 16'd44 )  ;
assign XRAM_addr_n1133 = n1132 ;
assign n1135 = XRAM_data_n1134 ;
assign n1136 =  { ( n1131 ) , ( n1135 ) }  ;
assign n1137 =  ( n912 ) + ( 16'd45 )  ;
assign XRAM_addr_n1138 = n1137 ;
assign n1140 = XRAM_data_n1139 ;
assign n1141 =  { ( n1136 ) , ( n1140 ) }  ;
assign n1142 =  ( n912 ) + ( 16'd46 )  ;
assign XRAM_addr_n1143 = n1142 ;
assign n1145 = XRAM_data_n1144 ;
assign n1146 =  { ( n1141 ) , ( n1145 ) }  ;
assign n1147 =  ( n912 ) + ( 16'd47 )  ;
assign XRAM_addr_n1148 = n1147 ;
assign n1150 = XRAM_data_n1149 ;
assign n1151 =  { ( n1146 ) , ( n1150 ) }  ;
assign n1152 =  ( n912 ) + ( 16'd48 )  ;
assign XRAM_addr_n1153 = n1152 ;
assign n1155 = XRAM_data_n1154 ;
assign n1156 =  { ( n1151 ) , ( n1155 ) }  ;
assign n1157 =  ( n912 ) + ( 16'd49 )  ;
assign XRAM_addr_n1158 = n1157 ;
assign n1160 = XRAM_data_n1159 ;
assign n1161 =  { ( n1156 ) , ( n1160 ) }  ;
assign n1162 =  ( n912 ) + ( 16'd50 )  ;
assign XRAM_addr_n1163 = n1162 ;
assign n1165 = XRAM_data_n1164 ;
assign n1166 =  { ( n1161 ) , ( n1165 ) }  ;
assign n1167 =  ( n912 ) + ( 16'd51 )  ;
assign XRAM_addr_n1168 = n1167 ;
assign n1170 = XRAM_data_n1169 ;
assign n1171 =  { ( n1166 ) , ( n1170 ) }  ;
assign n1172 =  ( n912 ) + ( 16'd52 )  ;
assign XRAM_addr_n1173 = n1172 ;
assign n1175 = XRAM_data_n1174 ;
assign n1176 =  { ( n1171 ) , ( n1175 ) }  ;
assign n1177 =  ( n912 ) + ( 16'd53 )  ;
assign XRAM_addr_n1178 = n1177 ;
assign n1180 = XRAM_data_n1179 ;
assign n1181 =  { ( n1176 ) , ( n1180 ) }  ;
assign n1182 =  ( n912 ) + ( 16'd54 )  ;
assign XRAM_addr_n1183 = n1182 ;
assign n1185 = XRAM_data_n1184 ;
assign n1186 =  { ( n1181 ) , ( n1185 ) }  ;
assign n1187 =  ( n912 ) + ( 16'd55 )  ;
assign XRAM_addr_n1188 = n1187 ;
assign n1190 = XRAM_data_n1189 ;
assign n1191 =  { ( n1186 ) , ( n1190 ) }  ;
assign n1192 =  ( n912 ) + ( 16'd56 )  ;
assign XRAM_addr_n1193 = n1192 ;
assign n1195 = XRAM_data_n1194 ;
assign n1196 =  { ( n1191 ) , ( n1195 ) }  ;
assign n1197 =  ( n912 ) + ( 16'd57 )  ;
assign XRAM_addr_n1198 = n1197 ;
assign n1200 = XRAM_data_n1199 ;
assign n1201 =  { ( n1196 ) , ( n1200 ) }  ;
assign n1202 =  ( n912 ) + ( 16'd58 )  ;
assign XRAM_addr_n1203 = n1202 ;
assign n1205 = XRAM_data_n1204 ;
assign n1206 =  { ( n1201 ) , ( n1205 ) }  ;
assign n1207 =  ( n912 ) + ( 16'd59 )  ;
assign XRAM_addr_n1208 = n1207 ;
assign n1210 = XRAM_data_n1209 ;
assign n1211 =  { ( n1206 ) , ( n1210 ) }  ;
assign n1212 =  ( n912 ) + ( 16'd60 )  ;
assign XRAM_addr_n1213 = n1212 ;
assign n1215 = XRAM_data_n1214 ;
assign n1216 =  { ( n1211 ) , ( n1215 ) }  ;
assign n1217 =  ( n912 ) + ( 16'd61 )  ;
assign XRAM_addr_n1218 = n1217 ;
assign n1220 = XRAM_data_n1219 ;
assign n1221 =  { ( n1216 ) , ( n1220 ) }  ;
assign n1222 =  ( n912 ) + ( 16'd62 )  ;
assign XRAM_addr_n1223 = n1222 ;
assign n1225 = XRAM_data_n1224 ;
assign n1226 =  { ( n1221 ) , ( n1225 ) }  ;
assign n1227 =  ( n912 ) + ( 16'd63 )  ;
assign XRAM_addr_n1228 = n1227 ;
assign n1230 = XRAM_data_n1229 ;
assign n1231 =  { ( n1226 ) , ( n1230 ) }  ;
assign n1232 =  ( n911 ) ? ( n1231 ) : ( sha_rd_data ) ;
assign n1233 = sha_rdaddr[15:8] ;
assign n1234 =  { ( n1233 ) , ( cmddata ) }  ;
assign n1235 = sha_rdaddr[7:0] ;
assign n1236 =  { ( cmddata ) , ( n1235 ) }  ;
assign n1237 =  ( n11 ) & (n125 )  ;
assign n1238 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n1239 =  ( n1237 ) & (n1238 )  ;
assign n1240 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n1241 =  ( n1237 ) & (n1240 )  ;
assign n1242 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n1243 =  ( n1237 ) & (n1242 )  ;
assign n1244 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n1245 =  ( n1237 ) & (n1244 )  ;
assign n1246 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n1247 =  ( n1237 ) & (n1246 )  ;
assign n1248 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n1249 =  ( n1237 ) & (n1248 )  ;
assign n1250 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n1251 =  ( n1237 ) & (n1250 )  ;
assign n1252 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n1253 =  ( n1237 ) & (n1252 )  ;
assign n1254 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n1255 =  ( n1237 ) & (n1254 )  ;
assign n1256 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n1257 =  ( n1237 ) & (n1256 )  ;
assign n1258 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n1259 =  ( n1237 ) & (n1258 )  ;
assign n1260 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n1261 =  ( n1237 ) & (n1260 )  ;
assign n1262 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n1263 =  ( n1237 ) & (n1262 )  ;
assign n1264 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n1265 =  ( n1237 ) & (n1264 )  ;
assign n1266 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n1267 =  ( n1237 ) & (n1266 )  ;
assign n1268 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n1269 =  ( n1237 ) & (n1268 )  ;
assign n1270 =  ( n11 ) & (n1 )  ;
assign n1271 =  ( n1270 ) & (n1238 )  ;
assign n1272 =  ( n1270 ) & (n1240 )  ;
assign n1273 =  ( n1270 ) & (n1242 )  ;
assign n1274 =  ( n1270 ) & (n1244 )  ;
assign n1275 =  ( n1270 ) & (n1246 )  ;
assign n1276 =  ( n1270 ) & (n1248 )  ;
assign n1277 =  ( n1270 ) & (n1250 )  ;
assign n1278 =  ( n1270 ) & (n1252 )  ;
assign n1279 =  ( n1270 ) & (n1254 )  ;
assign n1280 =  ( n1270 ) & (n1256 )  ;
assign n1281 =  ( n1270 ) & (n1258 )  ;
assign n1282 =  ( n1270 ) & (n1260 )  ;
assign n1283 =  ( n1270 ) & (n1262 )  ;
assign n1284 =  ( n1270 ) & (n1264 )  ;
assign n1285 =  ( n1270 ) & (n1266 )  ;
assign n1286 =  ( n1270 ) & (n1268 )  ;
assign n1287 =  ( n1285 ) | ( n1286 )  ;
assign n1288 =  ( n1284 ) | ( n1287 )  ;
assign n1289 =  ( n1283 ) | ( n1288 )  ;
assign n1290 =  ( n1282 ) | ( n1289 )  ;
assign n1291 =  ( n1281 ) | ( n1290 )  ;
assign n1292 =  ( n1280 ) | ( n1291 )  ;
assign n1293 =  ( n1279 ) | ( n1292 )  ;
assign n1294 =  ( n1278 ) | ( n1293 )  ;
assign n1295 =  ( n1277 ) | ( n1294 )  ;
assign n1296 =  ( n1276 ) | ( n1295 )  ;
assign n1297 =  ( n1275 ) | ( n1296 )  ;
assign n1298 =  ( n1274 ) | ( n1297 )  ;
assign n1299 =  ( n1273 ) | ( n1298 )  ;
assign n1300 =  ( n1272 ) | ( n1299 )  ;
assign n1301 =  ( n1271 ) | ( n1300 )  ;
assign n1302 =  ( n1269 ) | ( n1301 )  ;
assign n1303 =  ( n1267 ) | ( n1302 )  ;
assign n1304 =  ( n1265 ) | ( n1303 )  ;
assign n1305 =  ( n1263 ) | ( n1304 )  ;
assign n1306 =  ( n1261 ) | ( n1305 )  ;
assign n1307 =  ( n1259 ) | ( n1306 )  ;
assign n1308 =  ( n1257 ) | ( n1307 )  ;
assign n1309 =  ( n1255 ) | ( n1308 )  ;
assign n1310 =  ( n1253 ) | ( n1309 )  ;
assign n1311 =  ( n1251 ) | ( n1310 )  ;
assign n1312 =  ( n1249 ) | ( n1311 )  ;
assign n1313 =  ( n1247 ) | ( n1312 )  ;
assign n1314 =  ( n1245 ) | ( n1313 )  ;
assign n1315 =  ( n1243 ) | ( n1314 )  ;
assign n1316 =  ( n1241 ) | ( n1315 )  ;
assign n1317 =  ( n1239 ) | ( n1316 )  ;
assign n1318 =  ( sha_bytes_read ) < ( sha_len )  ;
assign n1319 =  ( n1318 ) ? ( 3'd1 ) : ( 3'd4 ) ;
assign n1320 =  ( n8 ) & (n125 )  ;
assign n1321 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n1322 =  ( n1320 ) & (n1321 )  ;
assign n1323 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n1324 =  ( n1320 ) & (n1323 )  ;
assign n1325 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n1326 =  ( n1320 ) & (n1325 )  ;
assign n1327 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n1328 =  ( n1320 ) & (n1327 )  ;
assign n1329 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n1330 =  ( n1320 ) & (n1329 )  ;
assign n1331 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n1332 =  ( n1320 ) & (n1331 )  ;
assign n1333 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n1334 =  ( n1320 ) & (n1333 )  ;
assign n1335 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n1336 =  ( n1320 ) & (n1335 )  ;
assign n1337 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n1338 =  ( n1320 ) & (n1337 )  ;
assign n1339 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n1340 =  ( n1320 ) & (n1339 )  ;
assign n1341 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n1342 =  ( n1320 ) & (n1341 )  ;
assign n1343 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n1344 =  ( n1320 ) & (n1343 )  ;
assign n1345 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n1346 =  ( n1320 ) & (n1345 )  ;
assign n1347 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n1348 =  ( n1320 ) & (n1347 )  ;
assign n1349 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n1350 =  ( n1320 ) & (n1349 )  ;
assign n1351 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n1352 =  ( n1320 ) & (n1351 )  ;
assign n1353 =  ( n8 ) & (n1 )  ;
assign n1354 =  ( n1353 ) & (n1321 )  ;
assign n1355 =  ( n1353 ) & (n1323 )  ;
assign n1356 =  ( n1353 ) & (n1325 )  ;
assign n1357 =  ( n1353 ) & (n1327 )  ;
assign n1358 =  ( n1353 ) & (n1329 )  ;
assign n1359 =  ( n1353 ) & (n1331 )  ;
assign n1360 =  ( n1353 ) & (n1333 )  ;
assign n1361 =  ( n1353 ) & (n1335 )  ;
assign n1362 =  ( n1353 ) & (n1337 )  ;
assign n1363 =  ( n1353 ) & (n1339 )  ;
assign n1364 =  ( n1353 ) & (n1341 )  ;
assign n1365 =  ( n1353 ) & (n1343 )  ;
assign n1366 =  ( n1353 ) & (n1345 )  ;
assign n1367 =  ( n1353 ) & (n1347 )  ;
assign n1368 =  ( n1353 ) & (n1349 )  ;
assign n1369 =  ( n1353 ) & (n1351 )  ;
assign n1370 =  ( n1368 ) | ( n1369 )  ;
assign n1371 =  ( n1367 ) | ( n1370 )  ;
assign n1372 =  ( n1366 ) | ( n1371 )  ;
assign n1373 =  ( n1365 ) | ( n1372 )  ;
assign n1374 =  ( n1364 ) | ( n1373 )  ;
assign n1375 =  ( n1363 ) | ( n1374 )  ;
assign n1376 =  ( n1362 ) | ( n1375 )  ;
assign n1377 =  ( n1361 ) | ( n1376 )  ;
assign n1378 =  ( n1360 ) | ( n1377 )  ;
assign n1379 =  ( n1359 ) | ( n1378 )  ;
assign n1380 =  ( n1358 ) | ( n1379 )  ;
assign n1381 =  ( n1357 ) | ( n1380 )  ;
assign n1382 =  ( n1356 ) | ( n1381 )  ;
assign n1383 =  ( n1355 ) | ( n1382 )  ;
assign n1384 =  ( n1354 ) | ( n1383 )  ;
assign n1385 =  ( n1352 ) | ( n1384 )  ;
assign n1386 =  ( n1350 ) | ( n1385 )  ;
assign n1387 =  ( n1348 ) | ( n1386 )  ;
assign n1388 =  ( n1346 ) | ( n1387 )  ;
assign n1389 =  ( n1344 ) | ( n1388 )  ;
assign n1390 =  ( n1342 ) | ( n1389 )  ;
assign n1391 =  ( n1340 ) | ( n1390 )  ;
assign n1392 =  ( n1338 ) | ( n1391 )  ;
assign n1393 =  ( n1336 ) | ( n1392 )  ;
assign n1394 =  ( n1334 ) | ( n1393 )  ;
assign n1395 =  ( n1332 ) | ( n1394 )  ;
assign n1396 =  ( n1330 ) | ( n1395 )  ;
assign n1397 =  ( n1328 ) | ( n1396 )  ;
assign n1398 =  ( n1326 ) | ( n1397 )  ;
assign n1399 =  ( n1324 ) | ( n1398 )  ;
assign n1400 =  ( n1322 ) | ( n1399 )  ;
assign n1401 =  ( n5 ) & (n125 )  ;
assign n1402 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n1403 =  ( n1401 ) & (n1402 )  ;
assign n1404 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n1405 =  ( n1401 ) & (n1404 )  ;
assign n1406 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n1407 =  ( n1401 ) & (n1406 )  ;
assign n1408 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n1409 =  ( n1401 ) & (n1408 )  ;
assign n1410 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n1411 =  ( n1401 ) & (n1410 )  ;
assign n1412 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n1413 =  ( n1401 ) & (n1412 )  ;
assign n1414 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n1415 =  ( n1401 ) & (n1414 )  ;
assign n1416 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n1417 =  ( n1401 ) & (n1416 )  ;
assign n1418 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n1419 =  ( n1401 ) & (n1418 )  ;
assign n1420 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n1421 =  ( n1401 ) & (n1420 )  ;
assign n1422 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n1423 =  ( n1401 ) & (n1422 )  ;
assign n1424 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n1425 =  ( n1401 ) & (n1424 )  ;
assign n1426 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n1427 =  ( n1401 ) & (n1426 )  ;
assign n1428 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n1429 =  ( n1401 ) & (n1428 )  ;
assign n1430 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n1431 =  ( n1401 ) & (n1430 )  ;
assign n1432 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n1433 =  ( n1401 ) & (n1432 )  ;
assign n1434 =  ( n5 ) & (n1 )  ;
assign n1435 =  ( n1434 ) & (n1402 )  ;
assign n1436 =  ( n1434 ) & (n1404 )  ;
assign n1437 =  ( n1434 ) & (n1406 )  ;
assign n1438 =  ( n1434 ) & (n1408 )  ;
assign n1439 =  ( n1434 ) & (n1410 )  ;
assign n1440 =  ( n1434 ) & (n1412 )  ;
assign n1441 =  ( n1434 ) & (n1414 )  ;
assign n1442 =  ( n1434 ) & (n1416 )  ;
assign n1443 =  ( n1434 ) & (n1418 )  ;
assign n1444 =  ( n1434 ) & (n1420 )  ;
assign n1445 =  ( n1434 ) & (n1422 )  ;
assign n1446 =  ( n1434 ) & (n1424 )  ;
assign n1447 =  ( n1434 ) & (n1426 )  ;
assign n1448 =  ( n1434 ) & (n1428 )  ;
assign n1449 =  ( n1434 ) & (n1430 )  ;
assign n1450 =  ( n1434 ) & (n1432 )  ;
assign n1451 =  ( n1449 ) | ( n1450 )  ;
assign n1452 =  ( n1448 ) | ( n1451 )  ;
assign n1453 =  ( n1447 ) | ( n1452 )  ;
assign n1454 =  ( n1446 ) | ( n1453 )  ;
assign n1455 =  ( n1445 ) | ( n1454 )  ;
assign n1456 =  ( n1444 ) | ( n1455 )  ;
assign n1457 =  ( n1443 ) | ( n1456 )  ;
assign n1458 =  ( n1442 ) | ( n1457 )  ;
assign n1459 =  ( n1441 ) | ( n1458 )  ;
assign n1460 =  ( n1440 ) | ( n1459 )  ;
assign n1461 =  ( n1439 ) | ( n1460 )  ;
assign n1462 =  ( n1438 ) | ( n1461 )  ;
assign n1463 =  ( n1437 ) | ( n1462 )  ;
assign n1464 =  ( n1436 ) | ( n1463 )  ;
assign n1465 =  ( n1435 ) | ( n1464 )  ;
assign n1466 =  ( n1433 ) | ( n1465 )  ;
assign n1467 =  ( n1431 ) | ( n1466 )  ;
assign n1468 =  ( n1429 ) | ( n1467 )  ;
assign n1469 =  ( n1427 ) | ( n1468 )  ;
assign n1470 =  ( n1425 ) | ( n1469 )  ;
assign n1471 =  ( n1423 ) | ( n1470 )  ;
assign n1472 =  ( n1421 ) | ( n1471 )  ;
assign n1473 =  ( n1419 ) | ( n1472 )  ;
assign n1474 =  ( n1417 ) | ( n1473 )  ;
assign n1475 =  ( n1415 ) | ( n1474 )  ;
assign n1476 =  ( n1413 ) | ( n1475 )  ;
assign n1477 =  ( n1411 ) | ( n1476 )  ;
assign n1478 =  ( n1409 ) | ( n1477 )  ;
assign n1479 =  ( n1407 ) | ( n1478 )  ;
assign n1480 =  ( n1405 ) | ( n1479 )  ;
assign n1481 =  ( n1403 ) | ( n1480 )  ;
assign n1482 =  ( sha_state ) == ( 3'd4 )  ;
assign n1483 = ~ ( n1 )  ;
assign n1484 =  ( n1482 ) & (n1483 )  ;
assign n1485 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n1486 =  ( n1484 ) & (n1485 )  ;
assign n1487 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n1488 =  ( n1484 ) & (n1487 )  ;
assign n1489 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n1490 =  ( n1484 ) & (n1489 )  ;
assign n1491 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n1492 =  ( n1484 ) & (n1491 )  ;
assign n1493 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n1494 =  ( n1484 ) & (n1493 )  ;
assign n1495 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n1496 =  ( n1484 ) & (n1495 )  ;
assign n1497 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n1498 =  ( n1484 ) & (n1497 )  ;
assign n1499 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n1500 =  ( n1484 ) & (n1499 )  ;
assign n1501 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n1502 =  ( n1484 ) & (n1501 )  ;
assign n1503 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n1504 =  ( n1484 ) & (n1503 )  ;
assign n1505 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n1506 =  ( n1484 ) & (n1505 )  ;
assign n1507 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n1508 =  ( n1484 ) & (n1507 )  ;
assign n1509 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n1510 =  ( n1484 ) & (n1509 )  ;
assign n1511 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n1512 =  ( n1484 ) & (n1511 )  ;
assign n1513 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n1514 =  ( n1484 ) & (n1513 )  ;
assign n1515 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n1516 =  ( n1484 ) & (n1515 )  ;
assign n1517 =  ( n0 ) & (n107 )  ;
assign n1518 =  ( n1517 ) & (n1485 )  ;
assign n1519 =  ( n1517 ) & (n1487 )  ;
assign n1520 =  ( n1517 ) & (n1489 )  ;
assign n1521 =  ( n1517 ) & (n1491 )  ;
assign n1522 =  ( n1517 ) & (n1493 )  ;
assign n1523 =  ( n1517 ) & (n1495 )  ;
assign n1524 =  ( n1517 ) & (n1497 )  ;
assign n1525 =  ( n1517 ) & (n1499 )  ;
assign n1526 =  ( n1517 ) & (n1501 )  ;
assign n1527 =  ( n1517 ) & (n1503 )  ;
assign n1528 =  ( n1517 ) & (n1505 )  ;
assign n1529 =  ( n1517 ) & (n1507 )  ;
assign n1530 =  ( n1517 ) & (n1509 )  ;
assign n1531 =  ( n1517 ) & (n1511 )  ;
assign n1532 =  ( n1517 ) & (n1513 )  ;
assign n1533 =  ( n1482 ) & (n738 )  ;
assign n1534 =  ( n1533 ) & (n1485 )  ;
assign n1535 =  ( n0 ) & (n1 )  ;
assign n1536 =  ( n1535 ) & (n1485 )  ;
assign n1537 =  ( n1533 ) & (n1487 )  ;
assign n1538 =  ( n1535 ) & (n1487 )  ;
assign n1539 =  ( n1533 ) & (n1489 )  ;
assign n1540 =  ( n1535 ) & (n1489 )  ;
assign n1541 =  ( n1533 ) & (n1491 )  ;
assign n1542 =  ( n1535 ) & (n1491 )  ;
assign n1543 =  ( n1533 ) & (n1493 )  ;
assign n1544 =  ( n1535 ) & (n1493 )  ;
assign n1545 =  ( n1533 ) & (n1495 )  ;
assign n1546 =  ( n1535 ) & (n1495 )  ;
assign n1547 =  ( n1533 ) & (n1497 )  ;
assign n1548 =  ( n1535 ) & (n1497 )  ;
assign n1549 =  ( n1533 ) & (n1499 )  ;
assign n1550 =  ( n1535 ) & (n1499 )  ;
assign n1551 =  ( n1533 ) & (n1501 )  ;
assign n1552 =  ( n1535 ) & (n1501 )  ;
assign n1553 =  ( n1533 ) & (n1503 )  ;
assign n1554 =  ( n1535 ) & (n1503 )  ;
assign n1555 =  ( n1533 ) & (n1505 )  ;
assign n1556 =  ( n1535 ) & (n1505 )  ;
assign n1557 =  ( n1533 ) & (n1507 )  ;
assign n1558 =  ( n1535 ) & (n1507 )  ;
assign n1559 =  ( n1533 ) & (n1509 )  ;
assign n1560 =  ( n1535 ) & (n1509 )  ;
assign n1561 =  ( n1533 ) & (n1511 )  ;
assign n1562 =  ( n1535 ) & (n1511 )  ;
assign n1563 =  ( n1533 ) & (n1513 )  ;
assign n1564 =  ( n1535 ) & (n1513 )  ;
assign n1565 =  ( n1533 ) & (n1515 )  ;
assign n1566 =  ( n1535 ) & (n1515 )  ;
assign n1567 =  ( n1565 ) | ( n1566 )  ;
assign n1568 =  ( n1564 ) | ( n1567 )  ;
assign n1569 =  ( n1563 ) | ( n1568 )  ;
assign n1570 =  ( n1562 ) | ( n1569 )  ;
assign n1571 =  ( n1561 ) | ( n1570 )  ;
assign n1572 =  ( n1560 ) | ( n1571 )  ;
assign n1573 =  ( n1559 ) | ( n1572 )  ;
assign n1574 =  ( n1558 ) | ( n1573 )  ;
assign n1575 =  ( n1557 ) | ( n1574 )  ;
assign n1576 =  ( n1556 ) | ( n1575 )  ;
assign n1577 =  ( n1555 ) | ( n1576 )  ;
assign n1578 =  ( n1554 ) | ( n1577 )  ;
assign n1579 =  ( n1553 ) | ( n1578 )  ;
assign n1580 =  ( n1552 ) | ( n1579 )  ;
assign n1581 =  ( n1551 ) | ( n1580 )  ;
assign n1582 =  ( n1550 ) | ( n1581 )  ;
assign n1583 =  ( n1549 ) | ( n1582 )  ;
assign n1584 =  ( n1548 ) | ( n1583 )  ;
assign n1585 =  ( n1547 ) | ( n1584 )  ;
assign n1586 =  ( n1546 ) | ( n1585 )  ;
assign n1587 =  ( n1545 ) | ( n1586 )  ;
assign n1588 =  ( n1544 ) | ( n1587 )  ;
assign n1589 =  ( n1543 ) | ( n1588 )  ;
assign n1590 =  ( n1542 ) | ( n1589 )  ;
assign n1591 =  ( n1541 ) | ( n1590 )  ;
assign n1592 =  ( n1540 ) | ( n1591 )  ;
assign n1593 =  ( n1539 ) | ( n1592 )  ;
assign n1594 =  ( n1538 ) | ( n1593 )  ;
assign n1595 =  ( n1537 ) | ( n1594 )  ;
assign n1596 =  ( n1536 ) | ( n1595 )  ;
assign n1597 =  ( n1534 ) | ( n1596 )  ;
assign n1598 =  ( n1532 ) | ( n1597 )  ;
assign n1599 =  ( n1531 ) | ( n1598 )  ;
assign n1600 =  ( n1530 ) | ( n1599 )  ;
assign n1601 =  ( n1529 ) | ( n1600 )  ;
assign n1602 =  ( n1528 ) | ( n1601 )  ;
assign n1603 =  ( n1527 ) | ( n1602 )  ;
assign n1604 =  ( n1526 ) | ( n1603 )  ;
assign n1605 =  ( n1525 ) | ( n1604 )  ;
assign n1606 =  ( n1524 ) | ( n1605 )  ;
assign n1607 =  ( n1523 ) | ( n1606 )  ;
assign n1608 =  ( n1522 ) | ( n1607 )  ;
assign n1609 =  ( n1521 ) | ( n1608 )  ;
assign n1610 =  ( n1520 ) | ( n1609 )  ;
assign n1611 =  ( n1519 ) | ( n1610 )  ;
assign n1612 =  ( n1518 ) | ( n1611 )  ;
assign n1613 =  ( n1516 ) | ( n1612 )  ;
assign n1614 =  ( n1514 ) | ( n1613 )  ;
assign n1615 =  ( n1512 ) | ( n1614 )  ;
assign n1616 =  ( n1510 ) | ( n1615 )  ;
assign n1617 =  ( n1508 ) | ( n1616 )  ;
assign n1618 =  ( n1506 ) | ( n1617 )  ;
assign n1619 =  ( n1504 ) | ( n1618 )  ;
assign n1620 =  ( n1502 ) | ( n1619 )  ;
assign n1621 =  ( n1500 ) | ( n1620 )  ;
assign n1622 =  ( n1498 ) | ( n1621 )  ;
assign n1623 =  ( n1496 ) | ( n1622 )  ;
assign n1624 =  ( n1494 ) | ( n1623 )  ;
assign n1625 =  ( n1492 ) | ( n1624 )  ;
assign n1626 =  ( n1490 ) | ( n1625 )  ;
assign n1627 =  ( n1488 ) | ( n1626 )  ;
assign n1628 =  ( n1486 ) | ( n1627 )  ;
assign n1629 =  ( n1628 ) ? ( 3'd0 ) : ( sha_state ) ;
assign n1630 =  ( n1481 ) ? ( 3'd2 ) : ( n1629 ) ;
assign n1631 =  ( n1400 ) ? ( 3'd3 ) : ( n1630 ) ;
assign n1632 =  ( n1317 ) ? ( n1319 ) : ( n1631 ) ;
assign n1633 =  ( cmddata ) == ( 8'd1 )  ;
assign n1634 =  ( n1633 ) ? ( 3'd1 ) : ( sha_state ) ;
assign n1635 = sha_wraddr[15:8] ;
assign n1636 =  { ( n1635 ) , ( cmddata ) }  ;
assign n1637 = sha_wraddr[7:0] ;
assign n1638 =  { ( cmddata ) , ( n1637 ) }  ;
assign n1639 = ~ ( n193 )  ;
assign n1640 =  ( 1'b1 ) & (n1639 )  ;
assign n1641 = ~ ( n192 )  ;
assign n1642 =  ( n1640 ) & (n1641 )  ;
assign n1643 = ~ ( n191 )  ;
assign n1644 =  ( n1642 ) & (n1643 )  ;
assign n1645 = ~ ( n190 )  ;
assign n1646 =  ( n1644 ) & (n1645 )  ;
assign n1647 = ~ ( n189 )  ;
assign n1648 =  ( n1646 ) & (n1647 )  ;
assign n1649 = ~ ( n188 )  ;
assign n1650 =  ( n1648 ) & (n1649 )  ;
assign n1651 = ~ ( n187 )  ;
assign n1652 =  ( n1650 ) & (n1651 )  ;
assign n1653 = ~ ( n186 )  ;
assign n1654 =  ( n1652 ) & (n1653 )  ;
assign n1655 = ~ ( n185 )  ;
assign n1656 =  ( n1654 ) & (n1655 )  ;
assign n1657 = ~ ( n184 )  ;
assign n1658 =  ( n1656 ) & (n1657 )  ;
assign n1659 = ~ ( n183 )  ;
assign n1660 =  ( n1658 ) & (n1659 )  ;
assign n1661 = ~ ( n182 )  ;
assign n1662 =  ( n1660 ) & (n1661 )  ;
assign n1663 = ~ ( n181 )  ;
assign n1664 =  ( n1662 ) & (n1663 )  ;
assign n1665 = ~ ( n180 )  ;
assign n1666 =  ( n1664 ) & (n1665 )  ;
assign n1667 = ~ ( n179 )  ;
assign n1668 =  ( n1666 ) & (n1667 )  ;
assign n1669 = ~ ( n178 )  ;
assign n1670 =  ( n1668 ) & (n1669 )  ;
assign n1671 = ~ ( n177 )  ;
assign n1672 =  ( n1670 ) & (n1671 )  ;
assign n1673 = ~ ( n176 )  ;
assign n1674 =  ( n1672 ) & (n1673 )  ;
assign n1675 = ~ ( n175 )  ;
assign n1676 =  ( n1674 ) & (n1675 )  ;
assign n1677 = ~ ( n174 )  ;
assign n1678 =  ( n1676 ) & (n1677 )  ;
assign n1679 = ~ ( n173 )  ;
assign n1680 =  ( n1678 ) & (n1679 )  ;
assign n1681 = ~ ( n172 )  ;
assign n1682 =  ( n1680 ) & (n1681 )  ;
assign n1683 = ~ ( n171 )  ;
assign n1684 =  ( n1682 ) & (n1683 )  ;
assign n1685 = ~ ( n170 )  ;
assign n1686 =  ( n1684 ) & (n1685 )  ;
assign n1687 = ~ ( n169 )  ;
assign n1688 =  ( n1686 ) & (n1687 )  ;
assign n1689 = ~ ( n168 )  ;
assign n1690 =  ( n1688 ) & (n1689 )  ;
assign n1691 = ~ ( n167 )  ;
assign n1692 =  ( n1690 ) & (n1691 )  ;
assign n1693 = ~ ( n166 )  ;
assign n1694 =  ( n1692 ) & (n1693 )  ;
assign n1695 = ~ ( n165 )  ;
assign n1696 =  ( n1694 ) & (n1695 )  ;
assign n1697 = ~ ( n164 )  ;
assign n1698 =  ( n1696 ) & (n1697 )  ;
assign n1699 = ~ ( n163 )  ;
assign n1700 =  ( n1698 ) & (n1699 )  ;
assign n1701 = ~ ( n162 )  ;
assign n1702 =  ( n1700 ) & (n1701 )  ;
assign n1703 = ~ ( n161 )  ;
assign n1704 =  ( n1702 ) & (n1703 )  ;
assign n1705 = ~ ( n160 )  ;
assign n1706 =  ( n1704 ) & (n1705 )  ;
assign n1707 = ~ ( n159 )  ;
assign n1708 =  ( n1706 ) & (n1707 )  ;
assign n1709 = ~ ( n158 )  ;
assign n1710 =  ( n1708 ) & (n1709 )  ;
assign n1711 = ~ ( n157 )  ;
assign n1712 =  ( n1710 ) & (n1711 )  ;
assign n1713 = ~ ( n156 )  ;
assign n1714 =  ( n1712 ) & (n1713 )  ;
assign n1715 = ~ ( n155 )  ;
assign n1716 =  ( n1714 ) & (n1715 )  ;
assign n1717 = ~ ( n154 )  ;
assign n1718 =  ( n1716 ) & (n1717 )  ;
assign n1719 = ~ ( n153 )  ;
assign n1720 =  ( n1718 ) & (n1719 )  ;
assign n1721 = ~ ( n152 )  ;
assign n1722 =  ( n1720 ) & (n1721 )  ;
assign n1723 = ~ ( n151 )  ;
assign n1724 =  ( n1722 ) & (n1723 )  ;
assign n1725 = ~ ( n150 )  ;
assign n1726 =  ( n1724 ) & (n1725 )  ;
assign n1727 = ~ ( n149 )  ;
assign n1728 =  ( n1726 ) & (n1727 )  ;
assign n1729 = ~ ( n148 )  ;
assign n1730 =  ( n1728 ) & (n1729 )  ;
assign n1731 = ~ ( n147 )  ;
assign n1732 =  ( n1730 ) & (n1731 )  ;
assign n1733 = ~ ( n146 )  ;
assign n1734 =  ( n1732 ) & (n1733 )  ;
assign n1735 = ~ ( n145 )  ;
assign n1736 =  ( n1734 ) & (n1735 )  ;
assign n1737 = ~ ( n144 )  ;
assign n1738 =  ( n1736 ) & (n1737 )  ;
assign n1739 = ~ ( n143 )  ;
assign n1740 =  ( n1738 ) & (n1739 )  ;
assign n1741 = ~ ( n142 )  ;
assign n1742 =  ( n1740 ) & (n1741 )  ;
assign n1743 = ~ ( n141 )  ;
assign n1744 =  ( n1742 ) & (n1743 )  ;
assign n1745 = ~ ( n140 )  ;
assign n1746 =  ( n1744 ) & (n1745 )  ;
assign n1747 = ~ ( n139 )  ;
assign n1748 =  ( n1746 ) & (n1747 )  ;
assign n1749 = ~ ( n138 )  ;
assign n1750 =  ( n1748 ) & (n1749 )  ;
assign n1751 = ~ ( n137 )  ;
assign n1752 =  ( n1750 ) & (n1751 )  ;
assign n1753 = ~ ( n136 )  ;
assign n1754 =  ( n1752 ) & (n1753 )  ;
assign n1755 = ~ ( n135 )  ;
assign n1756 =  ( n1754 ) & (n1755 )  ;
assign n1757 = ~ ( n134 )  ;
assign n1758 =  ( n1756 ) & (n1757 )  ;
assign n1759 = ~ ( n133 )  ;
assign n1760 =  ( n1758 ) & (n1759 )  ;
assign n1761 = ~ ( n131 )  ;
assign n1762 =  ( n1760 ) & (n1761 )  ;
assign n1763 = ~ ( n129 )  ;
assign n1764 =  ( n1762 ) & (n1763 )  ;
assign n1765 = ~ ( n127 )  ;
assign n1766 =  ( n1764 ) & (n1765 )  ;
assign n1767 = ~ ( n124 )  ;
assign n1768 =  ( n1766 ) & (n1767 )  ;
assign n1769 = ~ ( n123 )  ;
assign n1770 =  ( n1768 ) & (n1769 )  ;
assign n1771 = ~ ( n122 )  ;
assign n1772 =  ( n1770 ) & (n1771 )  ;
assign n1773 = ~ ( n121 )  ;
assign n1774 =  ( n1772 ) & (n1773 )  ;
assign n1775 = ~ ( n120 )  ;
assign n1776 =  ( n1774 ) & (n1775 )  ;
assign n1777 = ~ ( n119 )  ;
assign n1778 =  ( n1776 ) & (n1777 )  ;
assign n1779 = ~ ( n118 )  ;
assign n1780 =  ( n1778 ) & (n1779 )  ;
assign n1781 = ~ ( n117 )  ;
assign n1782 =  ( n1780 ) & (n1781 )  ;
assign n1783 = ~ ( n116 )  ;
assign n1784 =  ( n1782 ) & (n1783 )  ;
assign n1785 = ~ ( n115 )  ;
assign n1786 =  ( n1784 ) & (n1785 )  ;
assign n1787 = ~ ( n114 )  ;
assign n1788 =  ( n1786 ) & (n1787 )  ;
assign n1789 = ~ ( n113 )  ;
assign n1790 =  ( n1788 ) & (n1789 )  ;
assign n1791 = ~ ( n112 )  ;
assign n1792 =  ( n1790 ) & (n1791 )  ;
assign n1793 = ~ ( n111 )  ;
assign n1794 =  ( n1792 ) & (n1793 )  ;
assign n1795 = ~ ( n110 )  ;
assign n1796 =  ( n1794 ) & (n1795 )  ;
assign n1797 = ~ ( n109 )  ;
assign n1798 =  ( n1796 ) & (n1797 )  ;
assign n1799 = ~ ( n106 )  ;
assign n1800 =  ( n1798 ) & (n1799 )  ;
assign n1801 = ~ ( n105 )  ;
assign n1802 =  ( n1800 ) & (n1801 )  ;
assign n1803 = ~ ( n104 )  ;
assign n1804 =  ( n1802 ) & (n1803 )  ;
assign n1805 = ~ ( n103 )  ;
assign n1806 =  ( n1804 ) & (n1805 )  ;
assign n1807 = ~ ( n102 )  ;
assign n1808 =  ( n1806 ) & (n1807 )  ;
assign n1809 = ~ ( n100 )  ;
assign n1810 =  ( n1808 ) & (n1809 )  ;
assign n1811 = ~ ( n99 )  ;
assign n1812 =  ( n1810 ) & (n1811 )  ;
assign n1813 = ~ ( n98 )  ;
assign n1814 =  ( n1812 ) & (n1813 )  ;
assign n1815 = ~ ( n97 )  ;
assign n1816 =  ( n1814 ) & (n1815 )  ;
assign n1817 = ~ ( n96 )  ;
assign n1818 =  ( n1816 ) & (n1817 )  ;
assign n1819 = ~ ( n94 )  ;
assign n1820 =  ( n1818 ) & (n1819 )  ;
assign n1821 = ~ ( n93 )  ;
assign n1822 =  ( n1820 ) & (n1821 )  ;
assign n1823 = ~ ( n92 )  ;
assign n1824 =  ( n1822 ) & (n1823 )  ;
assign n1825 = ~ ( n91 )  ;
assign n1826 =  ( n1824 ) & (n1825 )  ;
assign n1827 = ~ ( n90 )  ;
assign n1828 =  ( n1826 ) & (n1827 )  ;
assign n1829 = ~ ( n88 )  ;
assign n1830 =  ( n1828 ) & (n1829 )  ;
assign n1831 = ~ ( n87 )  ;
assign n1832 =  ( n1830 ) & (n1831 )  ;
assign n1833 = ~ ( n86 )  ;
assign n1834 =  ( n1832 ) & (n1833 )  ;
assign n1835 = ~ ( n85 )  ;
assign n1836 =  ( n1834 ) & (n1835 )  ;
assign n1837 = ~ ( n84 )  ;
assign n1838 =  ( n1836 ) & (n1837 )  ;
assign n1839 = ~ ( n82 )  ;
assign n1840 =  ( n1838 ) & (n1839 )  ;
assign n1841 = ~ ( n81 )  ;
assign n1842 =  ( n1840 ) & (n1841 )  ;
assign n1843 = ~ ( n80 )  ;
assign n1844 =  ( n1842 ) & (n1843 )  ;
assign n1845 = ~ ( n79 )  ;
assign n1846 =  ( n1844 ) & (n1845 )  ;
assign n1847 = ~ ( n78 )  ;
assign n1848 =  ( n1846 ) & (n1847 )  ;
assign n1849 = ~ ( n76 )  ;
assign n1850 =  ( n1848 ) & (n1849 )  ;
assign n1851 = ~ ( n75 )  ;
assign n1852 =  ( n1850 ) & (n1851 )  ;
assign n1853 = ~ ( n74 )  ;
assign n1854 =  ( n1852 ) & (n1853 )  ;
assign n1855 = ~ ( n73 )  ;
assign n1856 =  ( n1854 ) & (n1855 )  ;
assign n1857 = ~ ( n72 )  ;
assign n1858 =  ( n1856 ) & (n1857 )  ;
assign n1859 = ~ ( n70 )  ;
assign n1860 =  ( n1858 ) & (n1859 )  ;
assign n1861 = ~ ( n69 )  ;
assign n1862 =  ( n1860 ) & (n1861 )  ;
assign n1863 = ~ ( n68 )  ;
assign n1864 =  ( n1862 ) & (n1863 )  ;
assign n1865 = ~ ( n67 )  ;
assign n1866 =  ( n1864 ) & (n1865 )  ;
assign n1867 = ~ ( n66 )  ;
assign n1868 =  ( n1866 ) & (n1867 )  ;
assign n1869 = ~ ( n64 )  ;
assign n1870 =  ( n1868 ) & (n1869 )  ;
assign n1871 = ~ ( n63 )  ;
assign n1872 =  ( n1870 ) & (n1871 )  ;
assign n1873 = ~ ( n62 )  ;
assign n1874 =  ( n1872 ) & (n1873 )  ;
assign n1875 = ~ ( n61 )  ;
assign n1876 =  ( n1874 ) & (n1875 )  ;
assign n1877 = ~ ( n60 )  ;
assign n1878 =  ( n1876 ) & (n1877 )  ;
assign n1879 = ~ ( n58 )  ;
assign n1880 =  ( n1878 ) & (n1879 )  ;
assign n1881 = ~ ( n57 )  ;
assign n1882 =  ( n1880 ) & (n1881 )  ;
assign n1883 = ~ ( n56 )  ;
assign n1884 =  ( n1882 ) & (n1883 )  ;
assign n1885 = ~ ( n55 )  ;
assign n1886 =  ( n1884 ) & (n1885 )  ;
assign n1887 = ~ ( n54 )  ;
assign n1888 =  ( n1886 ) & (n1887 )  ;
assign n1889 = ~ ( n52 )  ;
assign n1890 =  ( n1888 ) & (n1889 )  ;
assign n1891 = ~ ( n51 )  ;
assign n1892 =  ( n1890 ) & (n1891 )  ;
assign n1893 = ~ ( n50 )  ;
assign n1894 =  ( n1892 ) & (n1893 )  ;
assign n1895 = ~ ( n49 )  ;
assign n1896 =  ( n1894 ) & (n1895 )  ;
assign n1897 = ~ ( n48 )  ;
assign n1898 =  ( n1896 ) & (n1897 )  ;
assign n1899 = ~ ( n46 )  ;
assign n1900 =  ( n1898 ) & (n1899 )  ;
assign n1901 = ~ ( n45 )  ;
assign n1902 =  ( n1900 ) & (n1901 )  ;
assign n1903 = ~ ( n44 )  ;
assign n1904 =  ( n1902 ) & (n1903 )  ;
assign n1905 = ~ ( n43 )  ;
assign n1906 =  ( n1904 ) & (n1905 )  ;
assign n1907 = ~ ( n42 )  ;
assign n1908 =  ( n1906 ) & (n1907 )  ;
assign n1909 = ~ ( n40 )  ;
assign n1910 =  ( n1908 ) & (n1909 )  ;
assign n1911 = ~ ( n39 )  ;
assign n1912 =  ( n1910 ) & (n1911 )  ;
assign n1913 = ~ ( n38 )  ;
assign n1914 =  ( n1912 ) & (n1913 )  ;
assign n1915 = ~ ( n37 )  ;
assign n1916 =  ( n1914 ) & (n1915 )  ;
assign n1917 = ~ ( n36 )  ;
assign n1918 =  ( n1916 ) & (n1917 )  ;
assign n1919 = ~ ( n34 )  ;
assign n1920 =  ( n1918 ) & (n1919 )  ;
assign n1921 = ~ ( n33 )  ;
assign n1922 =  ( n1920 ) & (n1921 )  ;
assign n1923 = ~ ( n32 )  ;
assign n1924 =  ( n1922 ) & (n1923 )  ;
assign n1925 = ~ ( n31 )  ;
assign n1926 =  ( n1924 ) & (n1925 )  ;
assign n1927 = ~ ( n30 )  ;
assign n1928 =  ( n1926 ) & (n1927 )  ;
assign n1929 = ~ ( n28 )  ;
assign n1930 =  ( n1928 ) & (n1929 )  ;
assign n1931 = ~ ( n27 )  ;
assign n1932 =  ( n1930 ) & (n1931 )  ;
assign n1933 = ~ ( n26 )  ;
assign n1934 =  ( n1932 ) & (n1933 )  ;
assign n1935 = ~ ( n25 )  ;
assign n1936 =  ( n1934 ) & (n1935 )  ;
assign n1937 = ~ ( n24 )  ;
assign n1938 =  ( n1936 ) & (n1937 )  ;
assign n1939 = ~ ( n22 )  ;
assign n1940 =  ( n1938 ) & (n1939 )  ;
assign n1941 = ~ ( n21 )  ;
assign n1942 =  ( n1940 ) & (n1941 )  ;
assign n1943 = ~ ( n20 )  ;
assign n1944 =  ( n1942 ) & (n1943 )  ;
assign n1945 = ~ ( n19 )  ;
assign n1946 =  ( n1944 ) & (n1945 )  ;
assign n1947 = ~ ( n18 )  ;
assign n1948 =  ( n1946 ) & (n1947 )  ;
assign n1949 = ~ ( n16 )  ;
assign n1950 =  ( n1948 ) & (n1949 )  ;
assign n1951 = ~ ( n13 )  ;
assign n1952 =  ( n1950 ) & (n1951 )  ;
assign n1953 = ~ ( n10 )  ;
assign n1954 =  ( n1952 ) & (n1953 )  ;
assign n1955 = ~ ( n7 )  ;
assign n1956 =  ( n1954 ) & (n1955 )  ;
assign n1957 = ~ ( n4 )  ;
assign n1958 =  ( n1956 ) & (n1957 )  ;
assign n1959 =  ( n1956 ) & (n4 )  ;
assign n1960 =  ( n132 ) & (n101 )  ;
assign n1961 =  ( n130 ) & (n101 )  ;
assign n1962 =  ( n128 ) & (n101 )  ;
assign n1963 =  ( n126 ) & (n101 )  ;
assign n1964 =  ( n132 ) & (n95 )  ;
assign n1965 =  ( n130 ) & (n95 )  ;
assign n1966 =  ( n128 ) & (n95 )  ;
assign n1967 =  ( n126 ) & (n95 )  ;
assign n1968 =  ( n132 ) & (n89 )  ;
assign n1969 =  ( n130 ) & (n89 )  ;
assign n1970 =  ( n128 ) & (n89 )  ;
assign n1971 =  ( n126 ) & (n89 )  ;
assign n1972 =  ( n132 ) & (n83 )  ;
assign n1973 =  ( n130 ) & (n83 )  ;
assign n1974 =  ( n128 ) & (n83 )  ;
assign n1975 =  ( n126 ) & (n83 )  ;
assign n1976 =  ( n132 ) & (n77 )  ;
assign n1977 =  ( n130 ) & (n77 )  ;
assign n1978 =  ( n128 ) & (n77 )  ;
assign n1979 =  ( n126 ) & (n77 )  ;
assign n1980 =  ( n132 ) & (n71 )  ;
assign n1981 =  ( n130 ) & (n71 )  ;
assign n1982 =  ( n128 ) & (n71 )  ;
assign n1983 =  ( n126 ) & (n71 )  ;
assign n1984 =  ( n132 ) & (n65 )  ;
assign n1985 =  ( n130 ) & (n65 )  ;
assign n1986 =  ( n128 ) & (n65 )  ;
assign n1987 =  ( n126 ) & (n65 )  ;
assign n1988 =  ( n132 ) & (n59 )  ;
assign n1989 =  ( n130 ) & (n59 )  ;
assign n1990 =  ( n128 ) & (n59 )  ;
assign n1991 =  ( n126 ) & (n59 )  ;
assign n1992 =  ( n132 ) & (n53 )  ;
assign n1993 =  ( n130 ) & (n53 )  ;
assign n1994 =  ( n128 ) & (n53 )  ;
assign n1995 =  ( n126 ) & (n53 )  ;
assign n1996 =  ( n132 ) & (n47 )  ;
assign n1997 =  ( n130 ) & (n47 )  ;
assign n1998 =  ( n128 ) & (n47 )  ;
assign n1999 =  ( n126 ) & (n47 )  ;
assign n2000 =  ( n132 ) & (n41 )  ;
assign n2001 =  ( n130 ) & (n41 )  ;
assign n2002 =  ( n128 ) & (n41 )  ;
assign n2003 =  ( n126 ) & (n41 )  ;
assign n2004 =  ( n132 ) & (n35 )  ;
assign n2005 =  ( n130 ) & (n35 )  ;
assign n2006 =  ( n128 ) & (n35 )  ;
assign n2007 =  ( n126 ) & (n35 )  ;
assign n2008 =  ( n132 ) & (n29 )  ;
assign n2009 =  ( n130 ) & (n29 )  ;
assign n2010 =  ( n128 ) & (n29 )  ;
assign n2011 =  ( n126 ) & (n29 )  ;
assign n2012 =  ( n132 ) & (n23 )  ;
assign n2013 =  ( n130 ) & (n23 )  ;
assign n2014 =  ( n128 ) & (n23 )  ;
assign n2015 =  ( n126 ) & (n23 )  ;
assign n2016 =  ( n132 ) & (n17 )  ;
assign n2017 =  ( n130 ) & (n17 )  ;
assign n2018 =  ( n128 ) & (n17 )  ;
assign n2019 =  ( n126 ) & (n17 )  ;
assign n2020 =  ( n132 ) & (n3 )  ;
assign n2021 =  ( n130 ) & (n3 )  ;
assign n2022 =  ( n128 ) & (n3 )  ;
assign n2023 =  ( n126 ) & (n3 )  ;
assign n2024 =  ( n108 ) & (n101 )  ;
assign n2025 =  ( n108 ) & (n95 )  ;
assign n2026 =  ( n108 ) & (n89 )  ;
assign n2027 =  ( n108 ) & (n83 )  ;
assign n2028 =  ( n108 ) & (n77 )  ;
assign n2029 =  ( n108 ) & (n71 )  ;
assign n2030 =  ( n108 ) & (n65 )  ;
assign n2031 =  ( n108 ) & (n59 )  ;
assign n2032 =  ( n108 ) & (n53 )  ;
assign n2033 =  ( n108 ) & (n47 )  ;
assign n2034 =  ( n108 ) & (n41 )  ;
assign n2035 =  ( n108 ) & (n35 )  ;
assign n2036 =  ( n108 ) & (n29 )  ;
assign n2037 =  ( n108 ) & (n23 )  ;
assign n2038 =  ( n108 ) & (n17 )  ;
assign n2039 =  ( n108 ) & (n3 )  ;
assign n2040 =  ( n15 ) & (n101 )  ;
assign n2041 =  ( n12 ) & (n101 )  ;
assign n2042 =  ( n9 ) & (n101 )  ;
assign n2043 =  ( n6 ) & (n101 )  ;
assign n2044 =  ( n2 ) & (n101 )  ;
assign n2045 =  ( n15 ) & (n95 )  ;
assign n2046 =  ( n12 ) & (n95 )  ;
assign n2047 =  ( n9 ) & (n95 )  ;
assign n2048 =  ( n6 ) & (n95 )  ;
assign n2049 =  ( n2 ) & (n95 )  ;
assign n2050 =  ( n15 ) & (n89 )  ;
assign n2051 =  ( n12 ) & (n89 )  ;
assign n2052 =  ( n9 ) & (n89 )  ;
assign n2053 =  ( n6 ) & (n89 )  ;
assign n2054 =  ( n2 ) & (n89 )  ;
assign n2055 =  ( n15 ) & (n83 )  ;
assign n2056 =  ( n12 ) & (n83 )  ;
assign n2057 =  ( n9 ) & (n83 )  ;
assign n2058 =  ( n6 ) & (n83 )  ;
assign n2059 =  ( n2 ) & (n83 )  ;
assign n2060 =  ( n15 ) & (n77 )  ;
assign n2061 =  ( n12 ) & (n77 )  ;
assign n2062 =  ( n9 ) & (n77 )  ;
assign n2063 =  ( n6 ) & (n77 )  ;
assign n2064 =  ( n2 ) & (n77 )  ;
assign n2065 =  ( n15 ) & (n71 )  ;
assign n2066 =  ( n12 ) & (n71 )  ;
assign n2067 =  ( n9 ) & (n71 )  ;
assign n2068 =  ( n6 ) & (n71 )  ;
assign n2069 =  ( n2 ) & (n71 )  ;
assign n2070 =  ( n15 ) & (n65 )  ;
assign n2071 =  ( n12 ) & (n65 )  ;
assign n2072 =  ( n9 ) & (n65 )  ;
assign n2073 =  ( n6 ) & (n65 )  ;
assign n2074 =  ( n2 ) & (n65 )  ;
assign n2075 =  ( n15 ) & (n59 )  ;
assign n2076 =  ( n12 ) & (n59 )  ;
assign n2077 =  ( n9 ) & (n59 )  ;
assign n2078 =  ( n6 ) & (n59 )  ;
assign n2079 =  ( n2 ) & (n59 )  ;
assign n2080 =  ( n15 ) & (n53 )  ;
assign n2081 =  ( n12 ) & (n53 )  ;
assign n2082 =  ( n9 ) & (n53 )  ;
assign n2083 =  ( n6 ) & (n53 )  ;
assign n2084 =  ( n2 ) & (n53 )  ;
assign n2085 =  ( n15 ) & (n47 )  ;
assign n2086 =  ( n12 ) & (n47 )  ;
assign n2087 =  ( n9 ) & (n47 )  ;
assign n2088 =  ( n6 ) & (n47 )  ;
assign n2089 =  ( n2 ) & (n47 )  ;
assign n2090 =  ( n15 ) & (n41 )  ;
assign n2091 =  ( n12 ) & (n41 )  ;
assign n2092 =  ( n9 ) & (n41 )  ;
assign n2093 =  ( n6 ) & (n41 )  ;
assign n2094 =  ( n2 ) & (n41 )  ;
assign n2095 =  ( n15 ) & (n35 )  ;
assign n2096 =  ( n12 ) & (n35 )  ;
assign n2097 =  ( n9 ) & (n35 )  ;
assign n2098 =  ( n6 ) & (n35 )  ;
assign n2099 =  ( n2 ) & (n35 )  ;
assign n2100 =  ( n15 ) & (n29 )  ;
assign n2101 =  ( n12 ) & (n29 )  ;
assign n2102 =  ( n9 ) & (n29 )  ;
assign n2103 =  ( n6 ) & (n29 )  ;
assign n2104 =  ( n2 ) & (n29 )  ;
assign n2105 =  ( n15 ) & (n23 )  ;
assign n2106 =  ( n12 ) & (n23 )  ;
assign n2107 =  ( n9 ) & (n23 )  ;
assign n2108 =  ( n6 ) & (n23 )  ;
assign n2109 =  ( n2 ) & (n23 )  ;
assign n2110 =  ( n15 ) & (n17 )  ;
assign n2111 =  ( n12 ) & (n17 )  ;
assign n2112 =  ( n9 ) & (n17 )  ;
assign n2113 =  ( n6 ) & (n17 )  ;
assign n2114 =  ( n2 ) & (n17 )  ;
assign n2115 =  ( n15 ) & (n3 )  ;
assign n2116 =  ( n12 ) & (n3 )  ;
assign n2117 =  ( n9 ) & (n3 )  ;
assign n2118 =  ( n6 ) & (n3 )  ;
assign n2119 =  ( n2 ) & (n3 )  ;
assign n2120 =  ( n2118 ) | ( n2119 )  ;
assign n2121 =  ( n2117 ) | ( n2120 )  ;
assign n2122 =  ( n2116 ) | ( n2121 )  ;
assign n2123 =  ( n2115 ) | ( n2122 )  ;
assign n2124 =  ( n2114 ) | ( n2123 )  ;
assign n2125 =  ( n2113 ) | ( n2124 )  ;
assign n2126 =  ( n2112 ) | ( n2125 )  ;
assign n2127 =  ( n2111 ) | ( n2126 )  ;
assign n2128 =  ( n2110 ) | ( n2127 )  ;
assign n2129 =  ( n2109 ) | ( n2128 )  ;
assign n2130 =  ( n2108 ) | ( n2129 )  ;
assign n2131 =  ( n2107 ) | ( n2130 )  ;
assign n2132 =  ( n2106 ) | ( n2131 )  ;
assign n2133 =  ( n2105 ) | ( n2132 )  ;
assign n2134 =  ( n2104 ) | ( n2133 )  ;
assign n2135 =  ( n2103 ) | ( n2134 )  ;
assign n2136 =  ( n2102 ) | ( n2135 )  ;
assign n2137 =  ( n2101 ) | ( n2136 )  ;
assign n2138 =  ( n2100 ) | ( n2137 )  ;
assign n2139 =  ( n2099 ) | ( n2138 )  ;
assign n2140 =  ( n2098 ) | ( n2139 )  ;
assign n2141 =  ( n2097 ) | ( n2140 )  ;
assign n2142 =  ( n2096 ) | ( n2141 )  ;
assign n2143 =  ( n2095 ) | ( n2142 )  ;
assign n2144 =  ( n2094 ) | ( n2143 )  ;
assign n2145 =  ( n2093 ) | ( n2144 )  ;
assign n2146 =  ( n2092 ) | ( n2145 )  ;
assign n2147 =  ( n2091 ) | ( n2146 )  ;
assign n2148 =  ( n2090 ) | ( n2147 )  ;
assign n2149 =  ( n2089 ) | ( n2148 )  ;
assign n2150 =  ( n2088 ) | ( n2149 )  ;
assign n2151 =  ( n2087 ) | ( n2150 )  ;
assign n2152 =  ( n2086 ) | ( n2151 )  ;
assign n2153 =  ( n2085 ) | ( n2152 )  ;
assign n2154 =  ( n2084 ) | ( n2153 )  ;
assign n2155 =  ( n2083 ) | ( n2154 )  ;
assign n2156 =  ( n2082 ) | ( n2155 )  ;
assign n2157 =  ( n2081 ) | ( n2156 )  ;
assign n2158 =  ( n2080 ) | ( n2157 )  ;
assign n2159 =  ( n2079 ) | ( n2158 )  ;
assign n2160 =  ( n2078 ) | ( n2159 )  ;
assign n2161 =  ( n2077 ) | ( n2160 )  ;
assign n2162 =  ( n2076 ) | ( n2161 )  ;
assign n2163 =  ( n2075 ) | ( n2162 )  ;
assign n2164 =  ( n2074 ) | ( n2163 )  ;
assign n2165 =  ( n2073 ) | ( n2164 )  ;
assign n2166 =  ( n2072 ) | ( n2165 )  ;
assign n2167 =  ( n2071 ) | ( n2166 )  ;
assign n2168 =  ( n2070 ) | ( n2167 )  ;
assign n2169 =  ( n2069 ) | ( n2168 )  ;
assign n2170 =  ( n2068 ) | ( n2169 )  ;
assign n2171 =  ( n2067 ) | ( n2170 )  ;
assign n2172 =  ( n2066 ) | ( n2171 )  ;
assign n2173 =  ( n2065 ) | ( n2172 )  ;
assign n2174 =  ( n2064 ) | ( n2173 )  ;
assign n2175 =  ( n2063 ) | ( n2174 )  ;
assign n2176 =  ( n2062 ) | ( n2175 )  ;
assign n2177 =  ( n2061 ) | ( n2176 )  ;
assign n2178 =  ( n2060 ) | ( n2177 )  ;
assign n2179 =  ( n2059 ) | ( n2178 )  ;
assign n2180 =  ( n2058 ) | ( n2179 )  ;
assign n2181 =  ( n2057 ) | ( n2180 )  ;
assign n2182 =  ( n2056 ) | ( n2181 )  ;
assign n2183 =  ( n2055 ) | ( n2182 )  ;
assign n2184 =  ( n2054 ) | ( n2183 )  ;
assign n2185 =  ( n2053 ) | ( n2184 )  ;
assign n2186 =  ( n2052 ) | ( n2185 )  ;
assign n2187 =  ( n2051 ) | ( n2186 )  ;
assign n2188 =  ( n2050 ) | ( n2187 )  ;
assign n2189 =  ( n2049 ) | ( n2188 )  ;
assign n2190 =  ( n2048 ) | ( n2189 )  ;
assign n2191 =  ( n2047 ) | ( n2190 )  ;
assign n2192 =  ( n2046 ) | ( n2191 )  ;
assign n2193 =  ( n2045 ) | ( n2192 )  ;
assign n2194 =  ( n2044 ) | ( n2193 )  ;
assign n2195 =  ( n2043 ) | ( n2194 )  ;
assign n2196 =  ( n2042 ) | ( n2195 )  ;
assign n2197 =  ( n2041 ) | ( n2196 )  ;
assign n2198 =  ( n2040 ) | ( n2197 )  ;
assign n2199 =  ( n2039 ) | ( n2198 )  ;
assign n2200 =  ( n2038 ) | ( n2199 )  ;
assign n2201 =  ( n2037 ) | ( n2200 )  ;
assign n2202 =  ( n2036 ) | ( n2201 )  ;
assign n2203 =  ( n2035 ) | ( n2202 )  ;
assign n2204 =  ( n2034 ) | ( n2203 )  ;
assign n2205 =  ( n2033 ) | ( n2204 )  ;
assign n2206 =  ( n2032 ) | ( n2205 )  ;
assign n2207 =  ( n2031 ) | ( n2206 )  ;
assign n2208 =  ( n2030 ) | ( n2207 )  ;
assign n2209 =  ( n2029 ) | ( n2208 )  ;
assign n2210 =  ( n2028 ) | ( n2209 )  ;
assign n2211 =  ( n2027 ) | ( n2210 )  ;
assign n2212 =  ( n2026 ) | ( n2211 )  ;
assign n2213 =  ( n2025 ) | ( n2212 )  ;
assign n2214 =  ( n2024 ) | ( n2213 )  ;
assign n2215 =  ( n2023 ) | ( n2214 )  ;
assign n2216 =  ( n2022 ) | ( n2215 )  ;
assign n2217 =  ( n2021 ) | ( n2216 )  ;
assign n2218 =  ( n2020 ) | ( n2217 )  ;
assign n2219 =  ( n2019 ) | ( n2218 )  ;
assign n2220 =  ( n2018 ) | ( n2219 )  ;
assign n2221 =  ( n2017 ) | ( n2220 )  ;
assign n2222 =  ( n2016 ) | ( n2221 )  ;
assign n2223 =  ( n2015 ) | ( n2222 )  ;
assign n2224 =  ( n2014 ) | ( n2223 )  ;
assign n2225 =  ( n2013 ) | ( n2224 )  ;
assign n2226 =  ( n2012 ) | ( n2225 )  ;
assign n2227 =  ( n2011 ) | ( n2226 )  ;
assign n2228 =  ( n2010 ) | ( n2227 )  ;
assign n2229 =  ( n2009 ) | ( n2228 )  ;
assign n2230 =  ( n2008 ) | ( n2229 )  ;
assign n2231 =  ( n2007 ) | ( n2230 )  ;
assign n2232 =  ( n2006 ) | ( n2231 )  ;
assign n2233 =  ( n2005 ) | ( n2232 )  ;
assign n2234 =  ( n2004 ) | ( n2233 )  ;
assign n2235 =  ( n2003 ) | ( n2234 )  ;
assign n2236 =  ( n2002 ) | ( n2235 )  ;
assign n2237 =  ( n2001 ) | ( n2236 )  ;
assign n2238 =  ( n2000 ) | ( n2237 )  ;
assign n2239 =  ( n1999 ) | ( n2238 )  ;
assign n2240 =  ( n1998 ) | ( n2239 )  ;
assign n2241 =  ( n1997 ) | ( n2240 )  ;
assign n2242 =  ( n1996 ) | ( n2241 )  ;
assign n2243 =  ( n1995 ) | ( n2242 )  ;
assign n2244 =  ( n1994 ) | ( n2243 )  ;
assign n2245 =  ( n1993 ) | ( n2244 )  ;
assign n2246 =  ( n1992 ) | ( n2245 )  ;
assign n2247 =  ( n1991 ) | ( n2246 )  ;
assign n2248 =  ( n1990 ) | ( n2247 )  ;
assign n2249 =  ( n1989 ) | ( n2248 )  ;
assign n2250 =  ( n1988 ) | ( n2249 )  ;
assign n2251 =  ( n1987 ) | ( n2250 )  ;
assign n2252 =  ( n1986 ) | ( n2251 )  ;
assign n2253 =  ( n1985 ) | ( n2252 )  ;
assign n2254 =  ( n1984 ) | ( n2253 )  ;
assign n2255 =  ( n1983 ) | ( n2254 )  ;
assign n2256 =  ( n1982 ) | ( n2255 )  ;
assign n2257 =  ( n1981 ) | ( n2256 )  ;
assign n2258 =  ( n1980 ) | ( n2257 )  ;
assign n2259 =  ( n1979 ) | ( n2258 )  ;
assign n2260 =  ( n1978 ) | ( n2259 )  ;
assign n2261 =  ( n1977 ) | ( n2260 )  ;
assign n2262 =  ( n1976 ) | ( n2261 )  ;
assign n2263 =  ( n1975 ) | ( n2262 )  ;
assign n2264 =  ( n1974 ) | ( n2263 )  ;
assign n2265 =  ( n1973 ) | ( n2264 )  ;
assign n2266 =  ( n1972 ) | ( n2265 )  ;
assign n2267 =  ( n1971 ) | ( n2266 )  ;
assign n2268 =  ( n1970 ) | ( n2267 )  ;
assign n2269 =  ( n1969 ) | ( n2268 )  ;
assign n2270 =  ( n1968 ) | ( n2269 )  ;
assign n2271 =  ( n1967 ) | ( n2270 )  ;
assign n2272 =  ( n1966 ) | ( n2271 )  ;
assign n2273 =  ( n1965 ) | ( n2272 )  ;
assign n2274 =  ( n1964 ) | ( n2273 )  ;
assign n2275 =  ( n1963 ) | ( n2274 )  ;
assign n2276 =  ( n1962 ) | ( n2275 )  ;
assign n2277 =  ( n1961 ) | ( n2276 )  ;
assign n2278 =  ( n1960 ) | ( n2277 )  ;
assign n2279 = ~ ( n2278 )  ;
assign n2280 =  ( n1959 ) & (n2279 )  ;
assign n2281 =  ( n1959 ) & (n2278 )  ;
assign n2282 =  ( n14 ) & (n125 )  ;
assign n2283 =  ( cmdaddr ) == ( 16'd65039 )  ;
assign n2284 =  ( n2282 ) & (n2283 )  ;
assign n2285 =  ( cmdaddr ) == ( 16'd65038 )  ;
assign n2286 =  ( n2282 ) & (n2285 )  ;
assign n2287 =  ( cmdaddr ) == ( 16'd65037 )  ;
assign n2288 =  ( n2282 ) & (n2287 )  ;
assign n2289 =  ( cmdaddr ) == ( 16'd65036 )  ;
assign n2290 =  ( n2282 ) & (n2289 )  ;
assign n2291 =  ( cmdaddr ) == ( 16'd65035 )  ;
assign n2292 =  ( n2282 ) & (n2291 )  ;
assign n2293 =  ( cmdaddr ) == ( 16'd65034 )  ;
assign n2294 =  ( n2282 ) & (n2293 )  ;
assign n2295 =  ( cmdaddr ) == ( 16'd65033 )  ;
assign n2296 =  ( n2282 ) & (n2295 )  ;
assign n2297 =  ( cmdaddr ) == ( 16'd65032 )  ;
assign n2298 =  ( n2282 ) & (n2297 )  ;
assign n2299 =  ( cmdaddr ) == ( 16'd65031 )  ;
assign n2300 =  ( n2282 ) & (n2299 )  ;
assign n2301 =  ( cmdaddr ) == ( 16'd65030 )  ;
assign n2302 =  ( n2282 ) & (n2301 )  ;
assign n2303 =  ( cmdaddr ) == ( 16'd65029 )  ;
assign n2304 =  ( n2282 ) & (n2303 )  ;
assign n2305 =  ( cmdaddr ) == ( 16'd65028 )  ;
assign n2306 =  ( n2282 ) & (n2305 )  ;
assign n2307 =  ( cmdaddr ) == ( 16'd65027 )  ;
assign n2308 =  ( n2282 ) & (n2307 )  ;
assign n2309 =  ( cmdaddr ) == ( 16'd65026 )  ;
assign n2310 =  ( n2282 ) & (n2309 )  ;
assign n2311 =  ( cmdaddr ) == ( 16'd65025 )  ;
assign n2312 =  ( n2282 ) & (n2311 )  ;
assign n2313 =  ( cmdaddr ) == ( 16'd65024 )  ;
assign n2314 =  ( n2282 ) & (n2313 )  ;
assign n2315 =  ( n14 ) & (n1 )  ;
assign n2316 =  ( n2315 ) & (n2283 )  ;
assign n2317 =  ( n2315 ) & (n2285 )  ;
assign n2318 =  ( n2315 ) & (n2287 )  ;
assign n2319 =  ( n2315 ) & (n2289 )  ;
assign n2320 =  ( n2315 ) & (n2291 )  ;
assign n2321 =  ( n2315 ) & (n2293 )  ;
assign n2322 =  ( n2315 ) & (n2295 )  ;
assign n2323 =  ( n2315 ) & (n2297 )  ;
assign n2324 =  ( n2315 ) & (n2299 )  ;
assign n2325 =  ( n2315 ) & (n2301 )  ;
assign n2326 =  ( n2315 ) & (n2303 )  ;
assign n2327 =  ( n2315 ) & (n2305 )  ;
assign n2328 =  ( n2315 ) & (n2307 )  ;
assign n2329 =  ( n2315 ) & (n2309 )  ;
assign n2330 =  ( n2315 ) & (n2311 )  ;
assign n2331 =  ( n2315 ) & (n2313 )  ;
assign n2332 =  ( n2330 ) | ( n2331 )  ;
assign n2333 =  ( n2329 ) | ( n2332 )  ;
assign n2334 =  ( n2328 ) | ( n2333 )  ;
assign n2335 =  ( n2327 ) | ( n2334 )  ;
assign n2336 =  ( n2326 ) | ( n2335 )  ;
assign n2337 =  ( n2325 ) | ( n2336 )  ;
assign n2338 =  ( n2324 ) | ( n2337 )  ;
assign n2339 =  ( n2323 ) | ( n2338 )  ;
assign n2340 =  ( n2322 ) | ( n2339 )  ;
assign n2341 =  ( n2321 ) | ( n2340 )  ;
assign n2342 =  ( n2320 ) | ( n2341 )  ;
assign n2343 =  ( n2319 ) | ( n2342 )  ;
assign n2344 =  ( n2318 ) | ( n2343 )  ;
assign n2345 =  ( n2317 ) | ( n2344 )  ;
assign n2346 =  ( n2316 ) | ( n2345 )  ;
assign n2347 =  ( n2314 ) | ( n2346 )  ;
assign n2348 =  ( n2312 ) | ( n2347 )  ;
assign n2349 =  ( n2310 ) | ( n2348 )  ;
assign n2350 =  ( n2308 ) | ( n2349 )  ;
assign n2351 =  ( n2306 ) | ( n2350 )  ;
assign n2352 =  ( n2304 ) | ( n2351 )  ;
assign n2353 =  ( n2302 ) | ( n2352 )  ;
assign n2354 =  ( n2300 ) | ( n2353 )  ;
assign n2355 =  ( n2298 ) | ( n2354 )  ;
assign n2356 =  ( n2296 ) | ( n2355 )  ;
assign n2357 =  ( n2294 ) | ( n2356 )  ;
assign n2358 =  ( n2292 ) | ( n2357 )  ;
assign n2359 =  ( n2290 ) | ( n2358 )  ;
assign n2360 =  ( n2288 ) | ( n2359 )  ;
assign n2361 =  ( n2286 ) | ( n2360 )  ;
assign n2362 =  ( n2284 ) | ( n2361 )  ;
assign n2363 = ~ ( n2362 )  ;
assign n2364 =  ( n2281 ) & (n2363 )  ;
assign n2365 =  ( n2281 ) & (n2362 )  ;
assign n2366 =  ( sha_wraddr ) + ( 16'd7 )  ;
assign n2367 = sha_hs_data[103:96] ;
assign n2368 =  ( sha_wraddr ) + ( 16'd6 )  ;
assign n2369 = sha_hs_data[111:104] ;
assign n2370 =  ( sha_wraddr ) + ( 16'd5 )  ;
assign n2371 = sha_hs_data[119:112] ;
assign n2372 =  ( sha_wraddr ) + ( 16'd4 )  ;
assign n2373 = sha_hs_data[127:120] ;
assign n2374 =  ( sha_wraddr ) + ( 16'd3 )  ;
assign n2375 = sha_hs_data[135:128] ;
assign n2376 =  ( sha_wraddr ) + ( 16'd2 )  ;
assign n2377 = sha_hs_data[143:136] ;
assign n2378 =  ( sha_wraddr ) + ( 16'd1 )  ;
assign n2379 = sha_hs_data[151:144] ;
assign n2380 =  ( sha_wraddr ) + ( 16'd0 )  ;
assign n2381 = sha_hs_data[159:152] ;
assign n2382 =  ( n1954 ) & (n7 )  ;
assign n2383 = ~ ( n2278 )  ;
assign n2384 =  ( n2382 ) & (n2383 )  ;
assign n2385 =  ( n2382 ) & (n2278 )  ;
assign n2386 = ~ ( n2362 )  ;
assign n2387 =  ( n2385 ) & (n2386 )  ;
assign n2388 =  ( n2385 ) & (n2362 )  ;
assign n2389 =  ( n1952 ) & (n10 )  ;
assign n2390 = ~ ( n2278 )  ;
assign n2391 =  ( n2389 ) & (n2390 )  ;
assign n2392 =  ( n2389 ) & (n2278 )  ;
assign n2393 = ~ ( n2362 )  ;
assign n2394 =  ( n2392 ) & (n2393 )  ;
assign n2395 =  ( n2392 ) & (n2362 )  ;
assign n2396 =  ( n1950 ) & (n13 )  ;
assign n2397 = ~ ( n2278 )  ;
assign n2398 =  ( n2396 ) & (n2397 )  ;
assign n2399 =  ( n2396 ) & (n2278 )  ;
assign n2400 = ~ ( n2362 )  ;
assign n2401 =  ( n2399 ) & (n2400 )  ;
assign n2402 =  ( n2399 ) & (n2362 )  ;
assign n2403 =  ( n1948 ) & (n16 )  ;
assign n2404 = ~ ( n2278 )  ;
assign n2405 =  ( n2403 ) & (n2404 )  ;
assign n2406 =  ( n2403 ) & (n2278 )  ;
assign n2407 = ~ ( n2362 )  ;
assign n2408 =  ( n2406 ) & (n2407 )  ;
assign n2409 =  ( n2406 ) & (n2362 )  ;
assign n2410 =  ( n1946 ) & (n18 )  ;
assign n2411 = ~ ( n2278 )  ;
assign n2412 =  ( n2410 ) & (n2411 )  ;
assign n2413 =  ( n2410 ) & (n2278 )  ;
assign n2414 = ~ ( n2362 )  ;
assign n2415 =  ( n2413 ) & (n2414 )  ;
assign n2416 =  ( n2413 ) & (n2362 )  ;
assign n2417 =  ( n1944 ) & (n19 )  ;
assign n2418 = ~ ( n2278 )  ;
assign n2419 =  ( n2417 ) & (n2418 )  ;
assign n2420 =  ( n2417 ) & (n2278 )  ;
assign n2421 = ~ ( n2362 )  ;
assign n2422 =  ( n2420 ) & (n2421 )  ;
assign n2423 =  ( n2420 ) & (n2362 )  ;
assign n2424 =  ( n1942 ) & (n20 )  ;
assign n2425 = ~ ( n2278 )  ;
assign n2426 =  ( n2424 ) & (n2425 )  ;
assign n2427 =  ( n2424 ) & (n2278 )  ;
assign n2428 = ~ ( n2362 )  ;
assign n2429 =  ( n2427 ) & (n2428 )  ;
assign n2430 =  ( n2427 ) & (n2362 )  ;
assign n2431 =  ( n1940 ) & (n21 )  ;
assign n2432 = ~ ( n2278 )  ;
assign n2433 =  ( n2431 ) & (n2432 )  ;
assign n2434 =  ( n2431 ) & (n2278 )  ;
assign n2435 = ~ ( n2362 )  ;
assign n2436 =  ( n2434 ) & (n2435 )  ;
assign n2437 =  ( n2434 ) & (n2362 )  ;
assign n2438 =  ( n1938 ) & (n22 )  ;
assign n2439 = ~ ( n2278 )  ;
assign n2440 =  ( n2438 ) & (n2439 )  ;
assign n2441 =  ( n2438 ) & (n2278 )  ;
assign n2442 = ~ ( n2362 )  ;
assign n2443 =  ( n2441 ) & (n2442 )  ;
assign n2444 =  ( n2441 ) & (n2362 )  ;
assign n2445 =  ( n1936 ) & (n24 )  ;
assign n2446 = ~ ( n2278 )  ;
assign n2447 =  ( n2445 ) & (n2446 )  ;
assign n2448 =  ( n2445 ) & (n2278 )  ;
assign n2449 = ~ ( n2362 )  ;
assign n2450 =  ( n2448 ) & (n2449 )  ;
assign n2451 =  ( n2448 ) & (n2362 )  ;
assign n2452 =  ( n1934 ) & (n25 )  ;
assign n2453 = ~ ( n2278 )  ;
assign n2454 =  ( n2452 ) & (n2453 )  ;
assign n2455 =  ( n2452 ) & (n2278 )  ;
assign n2456 = ~ ( n2362 )  ;
assign n2457 =  ( n2455 ) & (n2456 )  ;
assign n2458 =  ( n2455 ) & (n2362 )  ;
assign n2459 =  ( n1932 ) & (n26 )  ;
assign n2460 = ~ ( n2278 )  ;
assign n2461 =  ( n2459 ) & (n2460 )  ;
assign n2462 =  ( n2459 ) & (n2278 )  ;
assign n2463 = ~ ( n2362 )  ;
assign n2464 =  ( n2462 ) & (n2463 )  ;
assign n2465 =  ( n2462 ) & (n2362 )  ;
assign n2466 =  ( n1930 ) & (n27 )  ;
assign n2467 = ~ ( n2278 )  ;
assign n2468 =  ( n2466 ) & (n2467 )  ;
assign n2469 =  ( n2466 ) & (n2278 )  ;
assign n2470 = ~ ( n2362 )  ;
assign n2471 =  ( n2469 ) & (n2470 )  ;
assign n2472 =  ( n2469 ) & (n2362 )  ;
assign n2473 =  ( n1928 ) & (n28 )  ;
assign n2474 = ~ ( n2278 )  ;
assign n2475 =  ( n2473 ) & (n2474 )  ;
assign n2476 =  ( n2473 ) & (n2278 )  ;
assign n2477 = ~ ( n2362 )  ;
assign n2478 =  ( n2476 ) & (n2477 )  ;
assign n2479 =  ( n2476 ) & (n2362 )  ;
assign n2480 =  ( n1926 ) & (n30 )  ;
assign n2481 = ~ ( n2278 )  ;
assign n2482 =  ( n2480 ) & (n2481 )  ;
assign n2483 =  ( n2480 ) & (n2278 )  ;
assign n2484 = ~ ( n2362 )  ;
assign n2485 =  ( n2483 ) & (n2484 )  ;
assign n2486 =  ( n2483 ) & (n2362 )  ;
assign n2487 =  ( n1924 ) & (n31 )  ;
assign n2488 = ~ ( n2278 )  ;
assign n2489 =  ( n2487 ) & (n2488 )  ;
assign n2490 =  ( n2487 ) & (n2278 )  ;
assign n2491 = ~ ( n2362 )  ;
assign n2492 =  ( n2490 ) & (n2491 )  ;
assign n2493 =  ( n2490 ) & (n2362 )  ;
assign n2494 =  ( n1922 ) & (n32 )  ;
assign n2495 = ~ ( n2278 )  ;
assign n2496 =  ( n2494 ) & (n2495 )  ;
assign n2497 =  ( n2494 ) & (n2278 )  ;
assign n2498 = ~ ( n2362 )  ;
assign n2499 =  ( n2497 ) & (n2498 )  ;
assign n2500 =  ( n2497 ) & (n2362 )  ;
assign n2501 =  ( n1920 ) & (n33 )  ;
assign n2502 = ~ ( n2278 )  ;
assign n2503 =  ( n2501 ) & (n2502 )  ;
assign n2504 =  ( n2501 ) & (n2278 )  ;
assign n2505 = ~ ( n2362 )  ;
assign n2506 =  ( n2504 ) & (n2505 )  ;
assign n2507 =  ( n2504 ) & (n2362 )  ;
assign n2508 =  ( n1918 ) & (n34 )  ;
assign n2509 = ~ ( n2278 )  ;
assign n2510 =  ( n2508 ) & (n2509 )  ;
assign n2511 =  ( n2508 ) & (n2278 )  ;
assign n2512 = ~ ( n2362 )  ;
assign n2513 =  ( n2511 ) & (n2512 )  ;
assign n2514 =  ( n2511 ) & (n2362 )  ;
assign n2515 =  ( n1916 ) & (n36 )  ;
assign n2516 = ~ ( n2278 )  ;
assign n2517 =  ( n2515 ) & (n2516 )  ;
assign n2518 =  ( n2515 ) & (n2278 )  ;
assign n2519 = ~ ( n2362 )  ;
assign n2520 =  ( n2518 ) & (n2519 )  ;
assign n2521 =  ( n2518 ) & (n2362 )  ;
assign n2522 =  ( n1914 ) & (n37 )  ;
assign n2523 = ~ ( n2278 )  ;
assign n2524 =  ( n2522 ) & (n2523 )  ;
assign n2525 =  ( n2522 ) & (n2278 )  ;
assign n2526 = ~ ( n2362 )  ;
assign n2527 =  ( n2525 ) & (n2526 )  ;
assign n2528 =  ( n2525 ) & (n2362 )  ;
assign n2529 =  ( n1912 ) & (n38 )  ;
assign n2530 = ~ ( n2278 )  ;
assign n2531 =  ( n2529 ) & (n2530 )  ;
assign n2532 =  ( n2529 ) & (n2278 )  ;
assign n2533 = ~ ( n2362 )  ;
assign n2534 =  ( n2532 ) & (n2533 )  ;
assign n2535 =  ( n2532 ) & (n2362 )  ;
assign n2536 =  ( n1910 ) & (n39 )  ;
assign n2537 = ~ ( n2278 )  ;
assign n2538 =  ( n2536 ) & (n2537 )  ;
assign n2539 =  ( n2536 ) & (n2278 )  ;
assign n2540 = ~ ( n2362 )  ;
assign n2541 =  ( n2539 ) & (n2540 )  ;
assign n2542 =  ( n2539 ) & (n2362 )  ;
assign n2543 =  ( n1908 ) & (n40 )  ;
assign n2544 = ~ ( n2278 )  ;
assign n2545 =  ( n2543 ) & (n2544 )  ;
assign n2546 =  ( n2543 ) & (n2278 )  ;
assign n2547 = ~ ( n2362 )  ;
assign n2548 =  ( n2546 ) & (n2547 )  ;
assign n2549 =  ( n2546 ) & (n2362 )  ;
assign n2550 =  ( n1906 ) & (n42 )  ;
assign n2551 = ~ ( n2278 )  ;
assign n2552 =  ( n2550 ) & (n2551 )  ;
assign n2553 =  ( n2550 ) & (n2278 )  ;
assign n2554 = ~ ( n2362 )  ;
assign n2555 =  ( n2553 ) & (n2554 )  ;
assign n2556 =  ( n2553 ) & (n2362 )  ;
assign n2557 =  ( n1904 ) & (n43 )  ;
assign n2558 = ~ ( n2278 )  ;
assign n2559 =  ( n2557 ) & (n2558 )  ;
assign n2560 =  ( n2557 ) & (n2278 )  ;
assign n2561 = ~ ( n2362 )  ;
assign n2562 =  ( n2560 ) & (n2561 )  ;
assign n2563 =  ( n2560 ) & (n2362 )  ;
assign n2564 =  ( n1902 ) & (n44 )  ;
assign n2565 = ~ ( n2278 )  ;
assign n2566 =  ( n2564 ) & (n2565 )  ;
assign n2567 =  ( n2564 ) & (n2278 )  ;
assign n2568 = ~ ( n2362 )  ;
assign n2569 =  ( n2567 ) & (n2568 )  ;
assign n2570 =  ( n2567 ) & (n2362 )  ;
assign n2571 =  ( n1900 ) & (n45 )  ;
assign n2572 = ~ ( n2278 )  ;
assign n2573 =  ( n2571 ) & (n2572 )  ;
assign n2574 =  ( n2571 ) & (n2278 )  ;
assign n2575 = ~ ( n2362 )  ;
assign n2576 =  ( n2574 ) & (n2575 )  ;
assign n2577 =  ( n2574 ) & (n2362 )  ;
assign n2578 =  ( n1898 ) & (n46 )  ;
assign n2579 = ~ ( n2278 )  ;
assign n2580 =  ( n2578 ) & (n2579 )  ;
assign n2581 =  ( n2578 ) & (n2278 )  ;
assign n2582 = ~ ( n2362 )  ;
assign n2583 =  ( n2581 ) & (n2582 )  ;
assign n2584 =  ( n2581 ) & (n2362 )  ;
assign n2585 =  ( n1896 ) & (n48 )  ;
assign n2586 = ~ ( n2278 )  ;
assign n2587 =  ( n2585 ) & (n2586 )  ;
assign n2588 =  ( n2585 ) & (n2278 )  ;
assign n2589 = ~ ( n2362 )  ;
assign n2590 =  ( n2588 ) & (n2589 )  ;
assign n2591 =  ( n2588 ) & (n2362 )  ;
assign n2592 =  ( n1894 ) & (n49 )  ;
assign n2593 = ~ ( n2278 )  ;
assign n2594 =  ( n2592 ) & (n2593 )  ;
assign n2595 =  ( n2592 ) & (n2278 )  ;
assign n2596 = ~ ( n2362 )  ;
assign n2597 =  ( n2595 ) & (n2596 )  ;
assign n2598 =  ( n2595 ) & (n2362 )  ;
assign n2599 =  ( n1892 ) & (n50 )  ;
assign n2600 = ~ ( n2278 )  ;
assign n2601 =  ( n2599 ) & (n2600 )  ;
assign n2602 =  ( n2599 ) & (n2278 )  ;
assign n2603 = ~ ( n2362 )  ;
assign n2604 =  ( n2602 ) & (n2603 )  ;
assign n2605 =  ( n2602 ) & (n2362 )  ;
assign n2606 =  ( n1890 ) & (n51 )  ;
assign n2607 = ~ ( n2278 )  ;
assign n2608 =  ( n2606 ) & (n2607 )  ;
assign n2609 =  ( n2606 ) & (n2278 )  ;
assign n2610 = ~ ( n2362 )  ;
assign n2611 =  ( n2609 ) & (n2610 )  ;
assign n2612 =  ( n2609 ) & (n2362 )  ;
assign n2613 =  ( n1888 ) & (n52 )  ;
assign n2614 = ~ ( n2278 )  ;
assign n2615 =  ( n2613 ) & (n2614 )  ;
assign n2616 =  ( n2613 ) & (n2278 )  ;
assign n2617 = ~ ( n2362 )  ;
assign n2618 =  ( n2616 ) & (n2617 )  ;
assign n2619 =  ( n2616 ) & (n2362 )  ;
assign n2620 =  ( n1886 ) & (n54 )  ;
assign n2621 = ~ ( n2278 )  ;
assign n2622 =  ( n2620 ) & (n2621 )  ;
assign n2623 =  ( n2620 ) & (n2278 )  ;
assign n2624 = ~ ( n2362 )  ;
assign n2625 =  ( n2623 ) & (n2624 )  ;
assign n2626 =  ( n2623 ) & (n2362 )  ;
assign n2627 =  ( n1884 ) & (n55 )  ;
assign n2628 = ~ ( n2278 )  ;
assign n2629 =  ( n2627 ) & (n2628 )  ;
assign n2630 =  ( n2627 ) & (n2278 )  ;
assign n2631 = ~ ( n2362 )  ;
assign n2632 =  ( n2630 ) & (n2631 )  ;
assign n2633 =  ( n2630 ) & (n2362 )  ;
assign n2634 =  ( n1882 ) & (n56 )  ;
assign n2635 = ~ ( n2278 )  ;
assign n2636 =  ( n2634 ) & (n2635 )  ;
assign n2637 =  ( n2634 ) & (n2278 )  ;
assign n2638 = ~ ( n2362 )  ;
assign n2639 =  ( n2637 ) & (n2638 )  ;
assign n2640 =  ( n2637 ) & (n2362 )  ;
assign n2641 =  ( n1880 ) & (n57 )  ;
assign n2642 = ~ ( n2278 )  ;
assign n2643 =  ( n2641 ) & (n2642 )  ;
assign n2644 =  ( n2641 ) & (n2278 )  ;
assign n2645 = ~ ( n2362 )  ;
assign n2646 =  ( n2644 ) & (n2645 )  ;
assign n2647 =  ( n2644 ) & (n2362 )  ;
assign n2648 =  ( n1878 ) & (n58 )  ;
assign n2649 = ~ ( n2278 )  ;
assign n2650 =  ( n2648 ) & (n2649 )  ;
assign n2651 =  ( n2648 ) & (n2278 )  ;
assign n2652 = ~ ( n2362 )  ;
assign n2653 =  ( n2651 ) & (n2652 )  ;
assign n2654 =  ( n2651 ) & (n2362 )  ;
assign n2655 =  ( n1876 ) & (n60 )  ;
assign n2656 = ~ ( n2278 )  ;
assign n2657 =  ( n2655 ) & (n2656 )  ;
assign n2658 =  ( n2655 ) & (n2278 )  ;
assign n2659 = ~ ( n2362 )  ;
assign n2660 =  ( n2658 ) & (n2659 )  ;
assign n2661 =  ( n2658 ) & (n2362 )  ;
assign n2662 =  ( n1874 ) & (n61 )  ;
assign n2663 = ~ ( n2278 )  ;
assign n2664 =  ( n2662 ) & (n2663 )  ;
assign n2665 =  ( n2662 ) & (n2278 )  ;
assign n2666 = ~ ( n2362 )  ;
assign n2667 =  ( n2665 ) & (n2666 )  ;
assign n2668 =  ( n2665 ) & (n2362 )  ;
assign n2669 =  ( n1872 ) & (n62 )  ;
assign n2670 = ~ ( n2278 )  ;
assign n2671 =  ( n2669 ) & (n2670 )  ;
assign n2672 =  ( n2669 ) & (n2278 )  ;
assign n2673 = ~ ( n2362 )  ;
assign n2674 =  ( n2672 ) & (n2673 )  ;
assign n2675 =  ( n2672 ) & (n2362 )  ;
assign n2676 =  ( n1870 ) & (n63 )  ;
assign n2677 = ~ ( n2278 )  ;
assign n2678 =  ( n2676 ) & (n2677 )  ;
assign n2679 =  ( n2676 ) & (n2278 )  ;
assign n2680 = ~ ( n2362 )  ;
assign n2681 =  ( n2679 ) & (n2680 )  ;
assign n2682 =  ( n2679 ) & (n2362 )  ;
assign n2683 =  ( n1868 ) & (n64 )  ;
assign n2684 = ~ ( n2278 )  ;
assign n2685 =  ( n2683 ) & (n2684 )  ;
assign n2686 =  ( n2683 ) & (n2278 )  ;
assign n2687 = ~ ( n2362 )  ;
assign n2688 =  ( n2686 ) & (n2687 )  ;
assign n2689 =  ( n2686 ) & (n2362 )  ;
assign n2690 =  ( n1866 ) & (n66 )  ;
assign n2691 = ~ ( n2278 )  ;
assign n2692 =  ( n2690 ) & (n2691 )  ;
assign n2693 =  ( n2690 ) & (n2278 )  ;
assign n2694 = ~ ( n2362 )  ;
assign n2695 =  ( n2693 ) & (n2694 )  ;
assign n2696 =  ( n2693 ) & (n2362 )  ;
assign n2697 =  ( n1864 ) & (n67 )  ;
assign n2698 = ~ ( n2278 )  ;
assign n2699 =  ( n2697 ) & (n2698 )  ;
assign n2700 =  ( n2697 ) & (n2278 )  ;
assign n2701 = ~ ( n2362 )  ;
assign n2702 =  ( n2700 ) & (n2701 )  ;
assign n2703 =  ( n2700 ) & (n2362 )  ;
assign n2704 =  ( n1862 ) & (n68 )  ;
assign n2705 = ~ ( n2278 )  ;
assign n2706 =  ( n2704 ) & (n2705 )  ;
assign n2707 =  ( n2704 ) & (n2278 )  ;
assign n2708 = ~ ( n2362 )  ;
assign n2709 =  ( n2707 ) & (n2708 )  ;
assign n2710 =  ( n2707 ) & (n2362 )  ;
assign n2711 =  ( n1860 ) & (n69 )  ;
assign n2712 = ~ ( n2278 )  ;
assign n2713 =  ( n2711 ) & (n2712 )  ;
assign n2714 =  ( n2711 ) & (n2278 )  ;
assign n2715 = ~ ( n2362 )  ;
assign n2716 =  ( n2714 ) & (n2715 )  ;
assign n2717 =  ( n2714 ) & (n2362 )  ;
assign n2718 =  ( n1858 ) & (n70 )  ;
assign n2719 = ~ ( n2278 )  ;
assign n2720 =  ( n2718 ) & (n2719 )  ;
assign n2721 =  ( n2718 ) & (n2278 )  ;
assign n2722 = ~ ( n2362 )  ;
assign n2723 =  ( n2721 ) & (n2722 )  ;
assign n2724 =  ( n2721 ) & (n2362 )  ;
assign n2725 =  ( n1856 ) & (n72 )  ;
assign n2726 = ~ ( n2278 )  ;
assign n2727 =  ( n2725 ) & (n2726 )  ;
assign n2728 =  ( n2725 ) & (n2278 )  ;
assign n2729 = ~ ( n2362 )  ;
assign n2730 =  ( n2728 ) & (n2729 )  ;
assign n2731 =  ( n2728 ) & (n2362 )  ;
assign n2732 =  ( n1854 ) & (n73 )  ;
assign n2733 = ~ ( n2278 )  ;
assign n2734 =  ( n2732 ) & (n2733 )  ;
assign n2735 =  ( n2732 ) & (n2278 )  ;
assign n2736 = ~ ( n2362 )  ;
assign n2737 =  ( n2735 ) & (n2736 )  ;
assign n2738 =  ( n2735 ) & (n2362 )  ;
assign n2739 =  ( n1852 ) & (n74 )  ;
assign n2740 = ~ ( n2278 )  ;
assign n2741 =  ( n2739 ) & (n2740 )  ;
assign n2742 =  ( n2739 ) & (n2278 )  ;
assign n2743 = ~ ( n2362 )  ;
assign n2744 =  ( n2742 ) & (n2743 )  ;
assign n2745 =  ( n2742 ) & (n2362 )  ;
assign n2746 =  ( n1850 ) & (n75 )  ;
assign n2747 = ~ ( n2278 )  ;
assign n2748 =  ( n2746 ) & (n2747 )  ;
assign n2749 =  ( n2746 ) & (n2278 )  ;
assign n2750 = ~ ( n2362 )  ;
assign n2751 =  ( n2749 ) & (n2750 )  ;
assign n2752 =  ( n2749 ) & (n2362 )  ;
assign n2753 =  ( n1848 ) & (n76 )  ;
assign n2754 = ~ ( n2278 )  ;
assign n2755 =  ( n2753 ) & (n2754 )  ;
assign n2756 =  ( n2753 ) & (n2278 )  ;
assign n2757 = ~ ( n2362 )  ;
assign n2758 =  ( n2756 ) & (n2757 )  ;
assign n2759 =  ( n2756 ) & (n2362 )  ;
assign n2760 =  ( n1846 ) & (n78 )  ;
assign n2761 = ~ ( n2278 )  ;
assign n2762 =  ( n2760 ) & (n2761 )  ;
assign n2763 =  ( n2760 ) & (n2278 )  ;
assign n2764 = ~ ( n2362 )  ;
assign n2765 =  ( n2763 ) & (n2764 )  ;
assign n2766 =  ( n2763 ) & (n2362 )  ;
assign n2767 =  ( n1844 ) & (n79 )  ;
assign n2768 = ~ ( n2278 )  ;
assign n2769 =  ( n2767 ) & (n2768 )  ;
assign n2770 =  ( n2767 ) & (n2278 )  ;
assign n2771 = ~ ( n2362 )  ;
assign n2772 =  ( n2770 ) & (n2771 )  ;
assign n2773 =  ( n2770 ) & (n2362 )  ;
assign n2774 =  ( n1842 ) & (n80 )  ;
assign n2775 = ~ ( n2278 )  ;
assign n2776 =  ( n2774 ) & (n2775 )  ;
assign n2777 =  ( n2774 ) & (n2278 )  ;
assign n2778 = ~ ( n2362 )  ;
assign n2779 =  ( n2777 ) & (n2778 )  ;
assign n2780 =  ( n2777 ) & (n2362 )  ;
assign n2781 =  ( n1840 ) & (n81 )  ;
assign n2782 = ~ ( n2278 )  ;
assign n2783 =  ( n2781 ) & (n2782 )  ;
assign n2784 =  ( n2781 ) & (n2278 )  ;
assign n2785 = ~ ( n2362 )  ;
assign n2786 =  ( n2784 ) & (n2785 )  ;
assign n2787 =  ( n2784 ) & (n2362 )  ;
assign n2788 =  ( n1838 ) & (n82 )  ;
assign n2789 = ~ ( n2278 )  ;
assign n2790 =  ( n2788 ) & (n2789 )  ;
assign n2791 =  ( n2788 ) & (n2278 )  ;
assign n2792 = ~ ( n2362 )  ;
assign n2793 =  ( n2791 ) & (n2792 )  ;
assign n2794 =  ( n2791 ) & (n2362 )  ;
assign n2795 =  ( n1836 ) & (n84 )  ;
assign n2796 = ~ ( n2278 )  ;
assign n2797 =  ( n2795 ) & (n2796 )  ;
assign n2798 =  ( n2795 ) & (n2278 )  ;
assign n2799 = ~ ( n2362 )  ;
assign n2800 =  ( n2798 ) & (n2799 )  ;
assign n2801 =  ( n2798 ) & (n2362 )  ;
assign n2802 =  ( n1834 ) & (n85 )  ;
assign n2803 = ~ ( n2278 )  ;
assign n2804 =  ( n2802 ) & (n2803 )  ;
assign n2805 =  ( n2802 ) & (n2278 )  ;
assign n2806 = ~ ( n2362 )  ;
assign n2807 =  ( n2805 ) & (n2806 )  ;
assign n2808 =  ( n2805 ) & (n2362 )  ;
assign n2809 =  ( n1832 ) & (n86 )  ;
assign n2810 = ~ ( n2278 )  ;
assign n2811 =  ( n2809 ) & (n2810 )  ;
assign n2812 =  ( n2809 ) & (n2278 )  ;
assign n2813 = ~ ( n2362 )  ;
assign n2814 =  ( n2812 ) & (n2813 )  ;
assign n2815 =  ( n2812 ) & (n2362 )  ;
assign n2816 =  ( n1830 ) & (n87 )  ;
assign n2817 = ~ ( n2278 )  ;
assign n2818 =  ( n2816 ) & (n2817 )  ;
assign n2819 =  ( n2816 ) & (n2278 )  ;
assign n2820 = ~ ( n2362 )  ;
assign n2821 =  ( n2819 ) & (n2820 )  ;
assign n2822 =  ( n2819 ) & (n2362 )  ;
assign n2823 =  ( n1828 ) & (n88 )  ;
assign n2824 = ~ ( n2278 )  ;
assign n2825 =  ( n2823 ) & (n2824 )  ;
assign n2826 =  ( n2823 ) & (n2278 )  ;
assign n2827 = ~ ( n2362 )  ;
assign n2828 =  ( n2826 ) & (n2827 )  ;
assign n2829 =  ( n2826 ) & (n2362 )  ;
assign n2830 =  ( n1826 ) & (n90 )  ;
assign n2831 = ~ ( n2278 )  ;
assign n2832 =  ( n2830 ) & (n2831 )  ;
assign n2833 =  ( n2830 ) & (n2278 )  ;
assign n2834 = ~ ( n2362 )  ;
assign n2835 =  ( n2833 ) & (n2834 )  ;
assign n2836 =  ( n2833 ) & (n2362 )  ;
assign n2837 =  ( n1824 ) & (n91 )  ;
assign n2838 = ~ ( n2278 )  ;
assign n2839 =  ( n2837 ) & (n2838 )  ;
assign n2840 =  ( n2837 ) & (n2278 )  ;
assign n2841 = ~ ( n2362 )  ;
assign n2842 =  ( n2840 ) & (n2841 )  ;
assign n2843 =  ( n2840 ) & (n2362 )  ;
assign n2844 =  ( n1822 ) & (n92 )  ;
assign n2845 = ~ ( n2278 )  ;
assign n2846 =  ( n2844 ) & (n2845 )  ;
assign n2847 =  ( n2844 ) & (n2278 )  ;
assign n2848 = ~ ( n2362 )  ;
assign n2849 =  ( n2847 ) & (n2848 )  ;
assign n2850 =  ( n2847 ) & (n2362 )  ;
assign n2851 =  ( n1820 ) & (n93 )  ;
assign n2852 = ~ ( n2278 )  ;
assign n2853 =  ( n2851 ) & (n2852 )  ;
assign n2854 =  ( n2851 ) & (n2278 )  ;
assign n2855 = ~ ( n2362 )  ;
assign n2856 =  ( n2854 ) & (n2855 )  ;
assign n2857 =  ( n2854 ) & (n2362 )  ;
assign n2858 =  ( n1818 ) & (n94 )  ;
assign n2859 = ~ ( n2278 )  ;
assign n2860 =  ( n2858 ) & (n2859 )  ;
assign n2861 =  ( n2858 ) & (n2278 )  ;
assign n2862 = ~ ( n2362 )  ;
assign n2863 =  ( n2861 ) & (n2862 )  ;
assign n2864 =  ( n2861 ) & (n2362 )  ;
assign n2865 =  ( n1816 ) & (n96 )  ;
assign n2866 = ~ ( n2278 )  ;
assign n2867 =  ( n2865 ) & (n2866 )  ;
assign n2868 =  ( n2865 ) & (n2278 )  ;
assign n2869 = ~ ( n2362 )  ;
assign n2870 =  ( n2868 ) & (n2869 )  ;
assign n2871 =  ( n2868 ) & (n2362 )  ;
assign n2872 =  ( n1814 ) & (n97 )  ;
assign n2873 = ~ ( n2278 )  ;
assign n2874 =  ( n2872 ) & (n2873 )  ;
assign n2875 =  ( n2872 ) & (n2278 )  ;
assign n2876 = ~ ( n2362 )  ;
assign n2877 =  ( n2875 ) & (n2876 )  ;
assign n2878 =  ( n2875 ) & (n2362 )  ;
assign n2879 =  ( n1812 ) & (n98 )  ;
assign n2880 = ~ ( n2278 )  ;
assign n2881 =  ( n2879 ) & (n2880 )  ;
assign n2882 =  ( n2879 ) & (n2278 )  ;
assign n2883 = ~ ( n2362 )  ;
assign n2884 =  ( n2882 ) & (n2883 )  ;
assign n2885 =  ( n2882 ) & (n2362 )  ;
assign n2886 =  ( n1810 ) & (n99 )  ;
assign n2887 = ~ ( n2278 )  ;
assign n2888 =  ( n2886 ) & (n2887 )  ;
assign n2889 =  ( n2886 ) & (n2278 )  ;
assign n2890 = ~ ( n2362 )  ;
assign n2891 =  ( n2889 ) & (n2890 )  ;
assign n2892 =  ( n2889 ) & (n2362 )  ;
assign n2893 =  ( n1808 ) & (n100 )  ;
assign n2894 = ~ ( n2278 )  ;
assign n2895 =  ( n2893 ) & (n2894 )  ;
assign n2896 =  ( n2893 ) & (n2278 )  ;
assign n2897 = ~ ( n2362 )  ;
assign n2898 =  ( n2896 ) & (n2897 )  ;
assign n2899 =  ( n2896 ) & (n2362 )  ;
assign n2900 =  ( n1806 ) & (n102 )  ;
assign n2901 = ~ ( n2278 )  ;
assign n2902 =  ( n2900 ) & (n2901 )  ;
assign n2903 =  ( n2900 ) & (n2278 )  ;
assign n2904 = ~ ( n2362 )  ;
assign n2905 =  ( n2903 ) & (n2904 )  ;
assign n2906 =  ( n2903 ) & (n2362 )  ;
assign n2907 =  ( n1804 ) & (n103 )  ;
assign n2908 = ~ ( n2278 )  ;
assign n2909 =  ( n2907 ) & (n2908 )  ;
assign n2910 =  ( n2907 ) & (n2278 )  ;
assign n2911 = ~ ( n2362 )  ;
assign n2912 =  ( n2910 ) & (n2911 )  ;
assign n2913 =  ( n2910 ) & (n2362 )  ;
assign n2914 =  ( n1802 ) & (n104 )  ;
assign n2915 = ~ ( n2278 )  ;
assign n2916 =  ( n2914 ) & (n2915 )  ;
assign n2917 =  ( n2914 ) & (n2278 )  ;
assign n2918 = ~ ( n2362 )  ;
assign n2919 =  ( n2917 ) & (n2918 )  ;
assign n2920 =  ( n2917 ) & (n2362 )  ;
assign n2921 =  ( n1800 ) & (n105 )  ;
assign n2922 = ~ ( n2278 )  ;
assign n2923 =  ( n2921 ) & (n2922 )  ;
assign n2924 =  ( n2921 ) & (n2278 )  ;
assign n2925 = ~ ( n2362 )  ;
assign n2926 =  ( n2924 ) & (n2925 )  ;
assign n2927 =  ( n2924 ) & (n2362 )  ;
assign n2928 =  ( n1798 ) & (n106 )  ;
assign n2929 = ~ ( n2278 )  ;
assign n2930 =  ( n2928 ) & (n2929 )  ;
assign n2931 =  ( n2928 ) & (n2278 )  ;
assign n2932 = ~ ( n2362 )  ;
assign n2933 =  ( n2931 ) & (n2932 )  ;
assign n2934 =  ( n2931 ) & (n2362 )  ;
assign n2935 =  ( n1796 ) & (n109 )  ;
assign n2936 = ~ ( n2278 )  ;
assign n2937 =  ( n2935 ) & (n2936 )  ;
assign n2938 =  ( n2935 ) & (n2278 )  ;
assign n2939 = ~ ( n2362 )  ;
assign n2940 =  ( n2938 ) & (n2939 )  ;
assign n2941 =  ( n2938 ) & (n2362 )  ;
assign n2942 =  ( n1794 ) & (n110 )  ;
assign n2943 = ~ ( n2278 )  ;
assign n2944 =  ( n2942 ) & (n2943 )  ;
assign n2945 =  ( n2942 ) & (n2278 )  ;
assign n2946 = ~ ( n2362 )  ;
assign n2947 =  ( n2945 ) & (n2946 )  ;
assign n2948 =  ( n2945 ) & (n2362 )  ;
assign n2949 =  ( n1792 ) & (n111 )  ;
assign n2950 = ~ ( n2278 )  ;
assign n2951 =  ( n2949 ) & (n2950 )  ;
assign n2952 =  ( n2949 ) & (n2278 )  ;
assign n2953 = ~ ( n2362 )  ;
assign n2954 =  ( n2952 ) & (n2953 )  ;
assign n2955 =  ( n2952 ) & (n2362 )  ;
assign n2956 =  ( n1790 ) & (n112 )  ;
assign n2957 = ~ ( n2278 )  ;
assign n2958 =  ( n2956 ) & (n2957 )  ;
assign n2959 =  ( n2956 ) & (n2278 )  ;
assign n2960 = ~ ( n2362 )  ;
assign n2961 =  ( n2959 ) & (n2960 )  ;
assign n2962 =  ( n2959 ) & (n2362 )  ;
assign n2963 =  ( n1788 ) & (n113 )  ;
assign n2964 = ~ ( n2278 )  ;
assign n2965 =  ( n2963 ) & (n2964 )  ;
assign n2966 =  ( n2963 ) & (n2278 )  ;
assign n2967 = ~ ( n2362 )  ;
assign n2968 =  ( n2966 ) & (n2967 )  ;
assign n2969 =  ( n2966 ) & (n2362 )  ;
assign n2970 =  ( n1786 ) & (n114 )  ;
assign n2971 = ~ ( n2278 )  ;
assign n2972 =  ( n2970 ) & (n2971 )  ;
assign n2973 =  ( n2970 ) & (n2278 )  ;
assign n2974 = ~ ( n2362 )  ;
assign n2975 =  ( n2973 ) & (n2974 )  ;
assign n2976 =  ( n2973 ) & (n2362 )  ;
assign n2977 =  ( n1784 ) & (n115 )  ;
assign n2978 = ~ ( n2278 )  ;
assign n2979 =  ( n2977 ) & (n2978 )  ;
assign n2980 =  ( n2977 ) & (n2278 )  ;
assign n2981 = ~ ( n2362 )  ;
assign n2982 =  ( n2980 ) & (n2981 )  ;
assign n2983 =  ( n2980 ) & (n2362 )  ;
assign n2984 =  ( n1782 ) & (n116 )  ;
assign n2985 = ~ ( n2278 )  ;
assign n2986 =  ( n2984 ) & (n2985 )  ;
assign n2987 =  ( n2984 ) & (n2278 )  ;
assign n2988 = ~ ( n2362 )  ;
assign n2989 =  ( n2987 ) & (n2988 )  ;
assign n2990 =  ( n2987 ) & (n2362 )  ;
assign n2991 =  ( n1780 ) & (n117 )  ;
assign n2992 = ~ ( n2278 )  ;
assign n2993 =  ( n2991 ) & (n2992 )  ;
assign n2994 =  ( n2991 ) & (n2278 )  ;
assign n2995 = ~ ( n2362 )  ;
assign n2996 =  ( n2994 ) & (n2995 )  ;
assign n2997 =  ( n2994 ) & (n2362 )  ;
assign n2998 =  ( n1778 ) & (n118 )  ;
assign n2999 = ~ ( n2278 )  ;
assign n3000 =  ( n2998 ) & (n2999 )  ;
assign n3001 =  ( n2998 ) & (n2278 )  ;
assign n3002 = ~ ( n2362 )  ;
assign n3003 =  ( n3001 ) & (n3002 )  ;
assign n3004 =  ( n3001 ) & (n2362 )  ;
assign n3005 =  ( n1776 ) & (n119 )  ;
assign n3006 = ~ ( n2278 )  ;
assign n3007 =  ( n3005 ) & (n3006 )  ;
assign n3008 =  ( n3005 ) & (n2278 )  ;
assign n3009 = ~ ( n2362 )  ;
assign n3010 =  ( n3008 ) & (n3009 )  ;
assign n3011 =  ( n3008 ) & (n2362 )  ;
assign n3012 =  ( n1774 ) & (n120 )  ;
assign n3013 = ~ ( n2278 )  ;
assign n3014 =  ( n3012 ) & (n3013 )  ;
assign n3015 =  ( n3012 ) & (n2278 )  ;
assign n3016 = ~ ( n2362 )  ;
assign n3017 =  ( n3015 ) & (n3016 )  ;
assign n3018 =  ( n3015 ) & (n2362 )  ;
assign n3019 =  ( n1772 ) & (n121 )  ;
assign n3020 = ~ ( n2278 )  ;
assign n3021 =  ( n3019 ) & (n3020 )  ;
assign n3022 =  ( n3019 ) & (n2278 )  ;
assign n3023 = ~ ( n2362 )  ;
assign n3024 =  ( n3022 ) & (n3023 )  ;
assign n3025 =  ( n3022 ) & (n2362 )  ;
assign n3026 =  ( n1770 ) & (n122 )  ;
assign n3027 = ~ ( n2278 )  ;
assign n3028 =  ( n3026 ) & (n3027 )  ;
assign n3029 =  ( n3026 ) & (n2278 )  ;
assign n3030 = ~ ( n2362 )  ;
assign n3031 =  ( n3029 ) & (n3030 )  ;
assign n3032 =  ( n3029 ) & (n2362 )  ;
assign n3033 =  ( n1768 ) & (n123 )  ;
assign n3034 = ~ ( n2278 )  ;
assign n3035 =  ( n3033 ) & (n3034 )  ;
assign n3036 =  ( n3033 ) & (n2278 )  ;
assign n3037 = ~ ( n2362 )  ;
assign n3038 =  ( n3036 ) & (n3037 )  ;
assign n3039 =  ( n3036 ) & (n2362 )  ;
assign n3040 =  ( n1766 ) & (n124 )  ;
assign n3041 = ~ ( n2278 )  ;
assign n3042 =  ( n3040 ) & (n3041 )  ;
assign n3043 =  ( n3040 ) & (n2278 )  ;
assign n3044 = ~ ( n2362 )  ;
assign n3045 =  ( n3043 ) & (n3044 )  ;
assign n3046 =  ( n3043 ) & (n2362 )  ;
assign n3047 =  ( n1764 ) & (n127 )  ;
assign n3048 = ~ ( n2278 )  ;
assign n3049 =  ( n3047 ) & (n3048 )  ;
assign n3050 =  ( n3047 ) & (n2278 )  ;
assign n3051 = ~ ( n2362 )  ;
assign n3052 =  ( n3050 ) & (n3051 )  ;
assign n3053 =  ( n3050 ) & (n2362 )  ;
assign n3054 =  ( n1762 ) & (n129 )  ;
assign n3055 = ~ ( n2278 )  ;
assign n3056 =  ( n3054 ) & (n3055 )  ;
assign n3057 =  ( n3054 ) & (n2278 )  ;
assign n3058 = ~ ( n2362 )  ;
assign n3059 =  ( n3057 ) & (n3058 )  ;
assign n3060 =  ( n3057 ) & (n2362 )  ;
assign n3061 =  ( n1760 ) & (n131 )  ;
assign n3062 = ~ ( n2278 )  ;
assign n3063 =  ( n3061 ) & (n3062 )  ;
assign n3064 =  ( n3061 ) & (n2278 )  ;
assign n3065 = ~ ( n2362 )  ;
assign n3066 =  ( n3064 ) & (n3065 )  ;
assign n3067 =  ( n3064 ) & (n2362 )  ;
assign n3068 =  ( n1758 ) & (n133 )  ;
assign n3069 = ~ ( n2278 )  ;
assign n3070 =  ( n3068 ) & (n3069 )  ;
assign n3071 =  ( n3068 ) & (n2278 )  ;
assign n3072 = ~ ( n2362 )  ;
assign n3073 =  ( n3071 ) & (n3072 )  ;
assign n3074 =  ( n3071 ) & (n2362 )  ;
assign n3075 =  ( n1756 ) & (n134 )  ;
assign n3076 = ~ ( n2278 )  ;
assign n3077 =  ( n3075 ) & (n3076 )  ;
assign n3078 =  ( n3075 ) & (n2278 )  ;
assign n3079 = ~ ( n2362 )  ;
assign n3080 =  ( n3078 ) & (n3079 )  ;
assign n3081 =  ( n3078 ) & (n2362 )  ;
assign n3082 =  ( n1754 ) & (n135 )  ;
assign n3083 = ~ ( n2278 )  ;
assign n3084 =  ( n3082 ) & (n3083 )  ;
assign n3085 =  ( n3082 ) & (n2278 )  ;
assign n3086 = ~ ( n2362 )  ;
assign n3087 =  ( n3085 ) & (n3086 )  ;
assign n3088 =  ( n3085 ) & (n2362 )  ;
assign n3089 =  ( n1752 ) & (n136 )  ;
assign n3090 = ~ ( n2278 )  ;
assign n3091 =  ( n3089 ) & (n3090 )  ;
assign n3092 =  ( n3089 ) & (n2278 )  ;
assign n3093 = ~ ( n2362 )  ;
assign n3094 =  ( n3092 ) & (n3093 )  ;
assign n3095 =  ( n3092 ) & (n2362 )  ;
assign n3096 =  ( n1750 ) & (n137 )  ;
assign n3097 = ~ ( n2278 )  ;
assign n3098 =  ( n3096 ) & (n3097 )  ;
assign n3099 =  ( n3096 ) & (n2278 )  ;
assign n3100 = ~ ( n2362 )  ;
assign n3101 =  ( n3099 ) & (n3100 )  ;
assign n3102 =  ( n3099 ) & (n2362 )  ;
assign n3103 =  ( n1748 ) & (n138 )  ;
assign n3104 = ~ ( n2278 )  ;
assign n3105 =  ( n3103 ) & (n3104 )  ;
assign n3106 =  ( n3103 ) & (n2278 )  ;
assign n3107 = ~ ( n2362 )  ;
assign n3108 =  ( n3106 ) & (n3107 )  ;
assign n3109 =  ( n3106 ) & (n2362 )  ;
assign n3110 =  ( n1746 ) & (n139 )  ;
assign n3111 = ~ ( n2278 )  ;
assign n3112 =  ( n3110 ) & (n3111 )  ;
assign n3113 =  ( n3110 ) & (n2278 )  ;
assign n3114 = ~ ( n2362 )  ;
assign n3115 =  ( n3113 ) & (n3114 )  ;
assign n3116 =  ( n3113 ) & (n2362 )  ;
assign n3117 =  ( n1744 ) & (n140 )  ;
assign n3118 = ~ ( n2278 )  ;
assign n3119 =  ( n3117 ) & (n3118 )  ;
assign n3120 =  ( n3117 ) & (n2278 )  ;
assign n3121 = ~ ( n2362 )  ;
assign n3122 =  ( n3120 ) & (n3121 )  ;
assign n3123 =  ( n3120 ) & (n2362 )  ;
assign n3124 =  ( n1742 ) & (n141 )  ;
assign n3125 = ~ ( n2278 )  ;
assign n3126 =  ( n3124 ) & (n3125 )  ;
assign n3127 =  ( n3124 ) & (n2278 )  ;
assign n3128 = ~ ( n2362 )  ;
assign n3129 =  ( n3127 ) & (n3128 )  ;
assign n3130 =  ( n3127 ) & (n2362 )  ;
assign n3131 =  ( n1740 ) & (n142 )  ;
assign n3132 = ~ ( n2278 )  ;
assign n3133 =  ( n3131 ) & (n3132 )  ;
assign n3134 =  ( n3131 ) & (n2278 )  ;
assign n3135 = ~ ( n2362 )  ;
assign n3136 =  ( n3134 ) & (n3135 )  ;
assign n3137 =  ( n3134 ) & (n2362 )  ;
assign n3138 =  ( n1738 ) & (n143 )  ;
assign n3139 = ~ ( n2278 )  ;
assign n3140 =  ( n3138 ) & (n3139 )  ;
assign n3141 =  ( n3138 ) & (n2278 )  ;
assign n3142 = ~ ( n2362 )  ;
assign n3143 =  ( n3141 ) & (n3142 )  ;
assign n3144 =  ( n3141 ) & (n2362 )  ;
assign n3145 =  ( n1736 ) & (n144 )  ;
assign n3146 = ~ ( n2278 )  ;
assign n3147 =  ( n3145 ) & (n3146 )  ;
assign n3148 =  ( n3145 ) & (n2278 )  ;
assign n3149 = ~ ( n2362 )  ;
assign n3150 =  ( n3148 ) & (n3149 )  ;
assign n3151 =  ( n3148 ) & (n2362 )  ;
assign n3152 =  ( n1734 ) & (n145 )  ;
assign n3153 = ~ ( n2278 )  ;
assign n3154 =  ( n3152 ) & (n3153 )  ;
assign n3155 =  ( n3152 ) & (n2278 )  ;
assign n3156 = ~ ( n2362 )  ;
assign n3157 =  ( n3155 ) & (n3156 )  ;
assign n3158 =  ( n3155 ) & (n2362 )  ;
assign n3159 =  ( n1732 ) & (n146 )  ;
assign n3160 = ~ ( n2278 )  ;
assign n3161 =  ( n3159 ) & (n3160 )  ;
assign n3162 =  ( n3159 ) & (n2278 )  ;
assign n3163 = ~ ( n2362 )  ;
assign n3164 =  ( n3162 ) & (n3163 )  ;
assign n3165 =  ( n3162 ) & (n2362 )  ;
assign n3166 =  ( n1730 ) & (n147 )  ;
assign n3167 = ~ ( n2278 )  ;
assign n3168 =  ( n3166 ) & (n3167 )  ;
assign n3169 =  ( n3166 ) & (n2278 )  ;
assign n3170 = ~ ( n2362 )  ;
assign n3171 =  ( n3169 ) & (n3170 )  ;
assign n3172 =  ( n3169 ) & (n2362 )  ;
assign n3173 =  ( n1728 ) & (n148 )  ;
assign n3174 = ~ ( n2278 )  ;
assign n3175 =  ( n3173 ) & (n3174 )  ;
assign n3176 =  ( n3173 ) & (n2278 )  ;
assign n3177 = ~ ( n2362 )  ;
assign n3178 =  ( n3176 ) & (n3177 )  ;
assign n3179 =  ( n3176 ) & (n2362 )  ;
assign n3180 =  ( n1726 ) & (n149 )  ;
assign n3181 = ~ ( n2278 )  ;
assign n3182 =  ( n3180 ) & (n3181 )  ;
assign n3183 =  ( n3180 ) & (n2278 )  ;
assign n3184 = ~ ( n2362 )  ;
assign n3185 =  ( n3183 ) & (n3184 )  ;
assign n3186 =  ( n3183 ) & (n2362 )  ;
assign n3187 =  ( n1724 ) & (n150 )  ;
assign n3188 = ~ ( n2278 )  ;
assign n3189 =  ( n3187 ) & (n3188 )  ;
assign n3190 =  ( n3187 ) & (n2278 )  ;
assign n3191 = ~ ( n2362 )  ;
assign n3192 =  ( n3190 ) & (n3191 )  ;
assign n3193 =  ( n3190 ) & (n2362 )  ;
assign n3194 =  ( n1722 ) & (n151 )  ;
assign n3195 = ~ ( n2278 )  ;
assign n3196 =  ( n3194 ) & (n3195 )  ;
assign n3197 =  ( n3194 ) & (n2278 )  ;
assign n3198 = ~ ( n2362 )  ;
assign n3199 =  ( n3197 ) & (n3198 )  ;
assign n3200 =  ( n3197 ) & (n2362 )  ;
assign n3201 =  ( n1720 ) & (n152 )  ;
assign n3202 = ~ ( n2278 )  ;
assign n3203 =  ( n3201 ) & (n3202 )  ;
assign n3204 =  ( n3201 ) & (n2278 )  ;
assign n3205 = ~ ( n2362 )  ;
assign n3206 =  ( n3204 ) & (n3205 )  ;
assign n3207 =  ( n3204 ) & (n2362 )  ;
assign n3208 =  ( n1718 ) & (n153 )  ;
assign n3209 = ~ ( n2278 )  ;
assign n3210 =  ( n3208 ) & (n3209 )  ;
assign n3211 =  ( n3208 ) & (n2278 )  ;
assign n3212 = ~ ( n2362 )  ;
assign n3213 =  ( n3211 ) & (n3212 )  ;
assign n3214 =  ( n3211 ) & (n2362 )  ;
assign n3215 =  ( n1716 ) & (n154 )  ;
assign n3216 = ~ ( n2278 )  ;
assign n3217 =  ( n3215 ) & (n3216 )  ;
assign n3218 =  ( n3215 ) & (n2278 )  ;
assign n3219 = ~ ( n2362 )  ;
assign n3220 =  ( n3218 ) & (n3219 )  ;
assign n3221 =  ( n3218 ) & (n2362 )  ;
assign n3222 =  ( n1714 ) & (n155 )  ;
assign n3223 = ~ ( n2278 )  ;
assign n3224 =  ( n3222 ) & (n3223 )  ;
assign n3225 =  ( n3222 ) & (n2278 )  ;
assign n3226 = ~ ( n2362 )  ;
assign n3227 =  ( n3225 ) & (n3226 )  ;
assign n3228 =  ( n3225 ) & (n2362 )  ;
assign n3229 =  ( n1712 ) & (n156 )  ;
assign n3230 = ~ ( n2278 )  ;
assign n3231 =  ( n3229 ) & (n3230 )  ;
assign n3232 =  ( n3229 ) & (n2278 )  ;
assign n3233 = ~ ( n2362 )  ;
assign n3234 =  ( n3232 ) & (n3233 )  ;
assign n3235 =  ( n3232 ) & (n2362 )  ;
assign n3236 =  ( n1710 ) & (n157 )  ;
assign n3237 = ~ ( n2278 )  ;
assign n3238 =  ( n3236 ) & (n3237 )  ;
assign n3239 =  ( n3236 ) & (n2278 )  ;
assign n3240 = ~ ( n2362 )  ;
assign n3241 =  ( n3239 ) & (n3240 )  ;
assign n3242 =  ( n3239 ) & (n2362 )  ;
assign n3243 =  ( n1708 ) & (n158 )  ;
assign n3244 = ~ ( n2278 )  ;
assign n3245 =  ( n3243 ) & (n3244 )  ;
assign n3246 =  ( n3243 ) & (n2278 )  ;
assign n3247 = ~ ( n2362 )  ;
assign n3248 =  ( n3246 ) & (n3247 )  ;
assign n3249 =  ( n3246 ) & (n2362 )  ;
assign n3250 =  ( n1706 ) & (n159 )  ;
assign n3251 = ~ ( n2278 )  ;
assign n3252 =  ( n3250 ) & (n3251 )  ;
assign n3253 =  ( n3250 ) & (n2278 )  ;
assign n3254 = ~ ( n2362 )  ;
assign n3255 =  ( n3253 ) & (n3254 )  ;
assign n3256 =  ( n3253 ) & (n2362 )  ;
assign n3257 =  ( n1704 ) & (n160 )  ;
assign n3258 = ~ ( n2278 )  ;
assign n3259 =  ( n3257 ) & (n3258 )  ;
assign n3260 =  ( n3257 ) & (n2278 )  ;
assign n3261 = ~ ( n2362 )  ;
assign n3262 =  ( n3260 ) & (n3261 )  ;
assign n3263 =  ( n3260 ) & (n2362 )  ;
assign n3264 =  ( n1702 ) & (n161 )  ;
assign n3265 = ~ ( n2278 )  ;
assign n3266 =  ( n3264 ) & (n3265 )  ;
assign n3267 =  ( n3264 ) & (n2278 )  ;
assign n3268 = ~ ( n2362 )  ;
assign n3269 =  ( n3267 ) & (n3268 )  ;
assign n3270 =  ( n3267 ) & (n2362 )  ;
assign n3271 =  ( n1700 ) & (n162 )  ;
assign n3272 = ~ ( n2278 )  ;
assign n3273 =  ( n3271 ) & (n3272 )  ;
assign n3274 =  ( n3271 ) & (n2278 )  ;
assign n3275 = ~ ( n2362 )  ;
assign n3276 =  ( n3274 ) & (n3275 )  ;
assign n3277 =  ( n3274 ) & (n2362 )  ;
assign n3278 =  ( n1698 ) & (n163 )  ;
assign n3279 = ~ ( n2278 )  ;
assign n3280 =  ( n3278 ) & (n3279 )  ;
assign n3281 =  ( n3278 ) & (n2278 )  ;
assign n3282 = ~ ( n2362 )  ;
assign n3283 =  ( n3281 ) & (n3282 )  ;
assign n3284 =  ( n3281 ) & (n2362 )  ;
assign n3285 =  ( n1696 ) & (n164 )  ;
assign n3286 = ~ ( n2278 )  ;
assign n3287 =  ( n3285 ) & (n3286 )  ;
assign n3288 =  ( n3285 ) & (n2278 )  ;
assign n3289 = ~ ( n2362 )  ;
assign n3290 =  ( n3288 ) & (n3289 )  ;
assign n3291 =  ( n3288 ) & (n2362 )  ;
assign n3292 =  ( n1694 ) & (n165 )  ;
assign n3293 = ~ ( n2278 )  ;
assign n3294 =  ( n3292 ) & (n3293 )  ;
assign n3295 =  ( n3292 ) & (n2278 )  ;
assign n3296 = ~ ( n2362 )  ;
assign n3297 =  ( n3295 ) & (n3296 )  ;
assign n3298 =  ( n3295 ) & (n2362 )  ;
assign n3299 =  ( n1692 ) & (n166 )  ;
assign n3300 = ~ ( n2278 )  ;
assign n3301 =  ( n3299 ) & (n3300 )  ;
assign n3302 =  ( n3299 ) & (n2278 )  ;
assign n3303 = ~ ( n2362 )  ;
assign n3304 =  ( n3302 ) & (n3303 )  ;
assign n3305 =  ( n3302 ) & (n2362 )  ;
assign n3306 =  ( n1690 ) & (n167 )  ;
assign n3307 = ~ ( n2278 )  ;
assign n3308 =  ( n3306 ) & (n3307 )  ;
assign n3309 =  ( n3306 ) & (n2278 )  ;
assign n3310 = ~ ( n2362 )  ;
assign n3311 =  ( n3309 ) & (n3310 )  ;
assign n3312 =  ( n3309 ) & (n2362 )  ;
assign n3313 =  ( n1688 ) & (n168 )  ;
assign n3314 = ~ ( n2278 )  ;
assign n3315 =  ( n3313 ) & (n3314 )  ;
assign n3316 =  ( n3313 ) & (n2278 )  ;
assign n3317 = ~ ( n2362 )  ;
assign n3318 =  ( n3316 ) & (n3317 )  ;
assign n3319 =  ( n3316 ) & (n2362 )  ;
assign n3320 =  ( n1686 ) & (n169 )  ;
assign n3321 = ~ ( n2278 )  ;
assign n3322 =  ( n3320 ) & (n3321 )  ;
assign n3323 =  ( n3320 ) & (n2278 )  ;
assign n3324 = ~ ( n2362 )  ;
assign n3325 =  ( n3323 ) & (n3324 )  ;
assign n3326 =  ( n3323 ) & (n2362 )  ;
assign n3327 =  ( n1684 ) & (n170 )  ;
assign n3328 = ~ ( n2278 )  ;
assign n3329 =  ( n3327 ) & (n3328 )  ;
assign n3330 =  ( n3327 ) & (n2278 )  ;
assign n3331 = ~ ( n2362 )  ;
assign n3332 =  ( n3330 ) & (n3331 )  ;
assign n3333 =  ( n3330 ) & (n2362 )  ;
assign n3334 =  ( n1682 ) & (n171 )  ;
assign n3335 = ~ ( n2278 )  ;
assign n3336 =  ( n3334 ) & (n3335 )  ;
assign n3337 =  ( n3334 ) & (n2278 )  ;
assign n3338 = ~ ( n2362 )  ;
assign n3339 =  ( n3337 ) & (n3338 )  ;
assign n3340 =  ( n3337 ) & (n2362 )  ;
assign n3341 =  ( n1680 ) & (n172 )  ;
assign n3342 = ~ ( n2278 )  ;
assign n3343 =  ( n3341 ) & (n3342 )  ;
assign n3344 =  ( n3341 ) & (n2278 )  ;
assign n3345 = ~ ( n2362 )  ;
assign n3346 =  ( n3344 ) & (n3345 )  ;
assign n3347 =  ( n3344 ) & (n2362 )  ;
assign n3348 =  ( n1678 ) & (n173 )  ;
assign n3349 = ~ ( n2278 )  ;
assign n3350 =  ( n3348 ) & (n3349 )  ;
assign n3351 =  ( n3348 ) & (n2278 )  ;
assign n3352 = ~ ( n2362 )  ;
assign n3353 =  ( n3351 ) & (n3352 )  ;
assign n3354 =  ( n3351 ) & (n2362 )  ;
assign n3355 =  ( n1676 ) & (n174 )  ;
assign n3356 = ~ ( n2278 )  ;
assign n3357 =  ( n3355 ) & (n3356 )  ;
assign n3358 =  ( n3355 ) & (n2278 )  ;
assign n3359 = ~ ( n2362 )  ;
assign n3360 =  ( n3358 ) & (n3359 )  ;
assign n3361 =  ( n3358 ) & (n2362 )  ;
assign n3362 =  ( n1674 ) & (n175 )  ;
assign n3363 = ~ ( n2278 )  ;
assign n3364 =  ( n3362 ) & (n3363 )  ;
assign n3365 =  ( n3362 ) & (n2278 )  ;
assign n3366 = ~ ( n2362 )  ;
assign n3367 =  ( n3365 ) & (n3366 )  ;
assign n3368 =  ( n3365 ) & (n2362 )  ;
assign n3369 =  ( n1672 ) & (n176 )  ;
assign n3370 = ~ ( n2278 )  ;
assign n3371 =  ( n3369 ) & (n3370 )  ;
assign n3372 =  ( n3369 ) & (n2278 )  ;
assign n3373 = ~ ( n2362 )  ;
assign n3374 =  ( n3372 ) & (n3373 )  ;
assign n3375 =  ( n3372 ) & (n2362 )  ;
assign n3376 =  ( n1670 ) & (n177 )  ;
assign n3377 = ~ ( n2278 )  ;
assign n3378 =  ( n3376 ) & (n3377 )  ;
assign n3379 =  ( n3376 ) & (n2278 )  ;
assign n3380 = ~ ( n2362 )  ;
assign n3381 =  ( n3379 ) & (n3380 )  ;
assign n3382 =  ( n3379 ) & (n2362 )  ;
assign n3383 =  ( n1668 ) & (n178 )  ;
assign n3384 = ~ ( n2278 )  ;
assign n3385 =  ( n3383 ) & (n3384 )  ;
assign n3386 =  ( n3383 ) & (n2278 )  ;
assign n3387 = ~ ( n2362 )  ;
assign n3388 =  ( n3386 ) & (n3387 )  ;
assign n3389 =  ( n3386 ) & (n2362 )  ;
assign n3390 =  ( n1666 ) & (n179 )  ;
assign n3391 = ~ ( n2278 )  ;
assign n3392 =  ( n3390 ) & (n3391 )  ;
assign n3393 =  ( n3390 ) & (n2278 )  ;
assign n3394 = ~ ( n2362 )  ;
assign n3395 =  ( n3393 ) & (n3394 )  ;
assign n3396 =  ( n3393 ) & (n2362 )  ;
assign n3397 =  ( n1664 ) & (n180 )  ;
assign n3398 = ~ ( n2278 )  ;
assign n3399 =  ( n3397 ) & (n3398 )  ;
assign n3400 =  ( n3397 ) & (n2278 )  ;
assign n3401 = ~ ( n2362 )  ;
assign n3402 =  ( n3400 ) & (n3401 )  ;
assign n3403 =  ( n3400 ) & (n2362 )  ;
assign n3404 =  ( n1662 ) & (n181 )  ;
assign n3405 = ~ ( n2278 )  ;
assign n3406 =  ( n3404 ) & (n3405 )  ;
assign n3407 =  ( n3404 ) & (n2278 )  ;
assign n3408 = ~ ( n2362 )  ;
assign n3409 =  ( n3407 ) & (n3408 )  ;
assign n3410 =  ( n3407 ) & (n2362 )  ;
assign n3411 =  ( n1660 ) & (n182 )  ;
assign n3412 = ~ ( n2278 )  ;
assign n3413 =  ( n3411 ) & (n3412 )  ;
assign n3414 =  ( n3411 ) & (n2278 )  ;
assign n3415 = ~ ( n2362 )  ;
assign n3416 =  ( n3414 ) & (n3415 )  ;
assign n3417 =  ( n3414 ) & (n2362 )  ;
assign n3418 =  ( n1658 ) & (n183 )  ;
assign n3419 = ~ ( n2278 )  ;
assign n3420 =  ( n3418 ) & (n3419 )  ;
assign n3421 =  ( n3418 ) & (n2278 )  ;
assign n3422 = ~ ( n2362 )  ;
assign n3423 =  ( n3421 ) & (n3422 )  ;
assign n3424 =  ( n3421 ) & (n2362 )  ;
assign n3425 =  ( n1656 ) & (n184 )  ;
assign n3426 = ~ ( n2278 )  ;
assign n3427 =  ( n3425 ) & (n3426 )  ;
assign n3428 =  ( n3425 ) & (n2278 )  ;
assign n3429 = ~ ( n2362 )  ;
assign n3430 =  ( n3428 ) & (n3429 )  ;
assign n3431 =  ( n3428 ) & (n2362 )  ;
assign n3432 =  ( n1654 ) & (n185 )  ;
assign n3433 = ~ ( n2278 )  ;
assign n3434 =  ( n3432 ) & (n3433 )  ;
assign n3435 =  ( n3432 ) & (n2278 )  ;
assign n3436 = ~ ( n2362 )  ;
assign n3437 =  ( n3435 ) & (n3436 )  ;
assign n3438 =  ( n3435 ) & (n2362 )  ;
assign n3439 =  ( n1652 ) & (n186 )  ;
assign n3440 = ~ ( n2278 )  ;
assign n3441 =  ( n3439 ) & (n3440 )  ;
assign n3442 =  ( n3439 ) & (n2278 )  ;
assign n3443 = ~ ( n2362 )  ;
assign n3444 =  ( n3442 ) & (n3443 )  ;
assign n3445 =  ( n3442 ) & (n2362 )  ;
assign n3446 =  ( n1650 ) & (n187 )  ;
assign n3447 = ~ ( n2278 )  ;
assign n3448 =  ( n3446 ) & (n3447 )  ;
assign n3449 =  ( n3446 ) & (n2278 )  ;
assign n3450 = ~ ( n2362 )  ;
assign n3451 =  ( n3449 ) & (n3450 )  ;
assign n3452 =  ( n3449 ) & (n2362 )  ;
assign n3453 =  ( n1648 ) & (n188 )  ;
assign n3454 = ~ ( n2278 )  ;
assign n3455 =  ( n3453 ) & (n3454 )  ;
assign n3456 =  ( n3453 ) & (n2278 )  ;
assign n3457 = ~ ( n2362 )  ;
assign n3458 =  ( n3456 ) & (n3457 )  ;
assign n3459 =  ( n3456 ) & (n2362 )  ;
assign n3460 =  ( n1646 ) & (n189 )  ;
assign n3461 = ~ ( n2278 )  ;
assign n3462 =  ( n3460 ) & (n3461 )  ;
assign n3463 =  ( n3460 ) & (n2278 )  ;
assign n3464 = ~ ( n2362 )  ;
assign n3465 =  ( n3463 ) & (n3464 )  ;
assign n3466 =  ( n3463 ) & (n2362 )  ;
assign n3467 =  ( n1644 ) & (n190 )  ;
assign n3468 = ~ ( n2278 )  ;
assign n3469 =  ( n3467 ) & (n3468 )  ;
assign n3470 =  ( n3467 ) & (n2278 )  ;
assign n3471 = ~ ( n2362 )  ;
assign n3472 =  ( n3470 ) & (n3471 )  ;
assign n3473 =  ( n3470 ) & (n2362 )  ;
assign n3474 =  ( n1642 ) & (n191 )  ;
assign n3475 = ~ ( n2278 )  ;
assign n3476 =  ( n3474 ) & (n3475 )  ;
assign n3477 =  ( n3474 ) & (n2278 )  ;
assign n3478 = ~ ( n2362 )  ;
assign n3479 =  ( n3477 ) & (n3478 )  ;
assign n3480 =  ( n3477 ) & (n2362 )  ;
assign n3481 =  ( n1640 ) & (n192 )  ;
assign n3482 = ~ ( n2278 )  ;
assign n3483 =  ( n3481 ) & (n3482 )  ;
assign n3484 =  ( n3481 ) & (n2278 )  ;
assign n3485 = ~ ( n2362 )  ;
assign n3486 =  ( n3484 ) & (n3485 )  ;
assign n3487 =  ( n3484 ) & (n2362 )  ;
assign n3488 =  ( 1'b1 ) & (n193 )  ;
assign n3489 = ~ ( n2278 )  ;
assign n3490 =  ( n3488 ) & (n3489 )  ;
assign n3491 =  ( n3488 ) & (n2278 )  ;
assign n3492 = ~ ( n2362 )  ;
assign n3493 =  ( n3491 ) & (n3492 )  ;
assign n3494 =  ( n3491 ) & (n2362 )  ;
assign XRAM_addr0 = n3494 ? (n2366) : (n3487 ? (n2366) : (n3480 ? (n2366) : (n3473 ? (n2366) : (n3466 ? (n2366) : (n3459 ? (n2366) : (n3452 ? (n2366) : (n3445 ? (n2366) : (n3438 ? (n2366) : (n3431 ? (n2366) : (n3424 ? (n2366) : (n3417 ? (n2366) : (n3410 ? (n2366) : (n3403 ? (n2366) : (n3396 ? (n2366) : (n3389 ? (n2366) : (n3382 ? (n2366) : (n3375 ? (n2366) : (n3368 ? (n2366) : (n3361 ? (n2366) : (n3354 ? (n2366) : (n3347 ? (n2366) : (n3340 ? (n2366) : (n3333 ? (n2366) : (n3326 ? (n2366) : (n3319 ? (n2366) : (n3312 ? (n2366) : (n3305 ? (n2366) : (n3298 ? (n2366) : (n3291 ? (n2366) : (n3284 ? (n2366) : (n3277 ? (n2366) : (n3270 ? (n2366) : (n3263 ? (n2366) : (n3256 ? (n2366) : (n3249 ? (n2366) : (n3242 ? (n2366) : (n3235 ? (n2366) : (n3228 ? (n2366) : (n3221 ? (n2366) : (n3214 ? (n2366) : (n3207 ? (n2366) : (n3200 ? (n2366) : (n3193 ? (n2366) : (n3186 ? (n2366) : (n3179 ? (n2366) : (n3172 ? (n2366) : (n3165 ? (n2366) : (n3158 ? (n2366) : (n3151 ? (n2366) : (n3144 ? (n2366) : (n3137 ? (n2366) : (n3130 ? (n2366) : (n3123 ? (n2366) : (n3116 ? (n2366) : (n3109 ? (n2366) : (n3102 ? (n2366) : (n3095 ? (n2366) : (n3088 ? (n2366) : (n3081 ? (n2366) : (n3074 ? (n2366) : (n3067 ? (n2366) : (n3060 ? (n2366) : (n3053 ? (n2366) : (n3046 ? (n2366) : (n3039 ? (n2366) : (n3032 ? (n2366) : (n3025 ? (n2366) : (n3018 ? (n2366) : (n3011 ? (n2366) : (n3004 ? (n2366) : (n2997 ? (n2366) : (n2990 ? (n2366) : (n2983 ? (n2366) : (n2976 ? (n2366) : (n2969 ? (n2366) : (n2962 ? (n2366) : (n2955 ? (n2366) : (n2948 ? (n2366) : (n2941 ? (n2366) : (n2934 ? (n2366) : (n2927 ? (n2366) : (n2920 ? (n2366) : (n2913 ? (n2366) : (n2906 ? (n2366) : (n2899 ? (n2366) : (n2892 ? (n2366) : (n2885 ? (n2366) : (n2878 ? (n2366) : (n2871 ? (n2366) : (n2864 ? (n2366) : (n2857 ? (n2366) : (n2850 ? (n2366) : (n2843 ? (n2366) : (n2836 ? (n2366) : (n2829 ? (n2366) : (n2822 ? (n2366) : (n2815 ? (n2366) : (n2808 ? (n2366) : (n2801 ? (n2366) : (n2794 ? (n2366) : (n2787 ? (n2366) : (n2780 ? (n2366) : (n2773 ? (n2366) : (n2766 ? (n2366) : (n2759 ? (n2366) : (n2752 ? (n2366) : (n2745 ? (n2366) : (n2738 ? (n2366) : (n2731 ? (n2366) : (n2724 ? (n2366) : (n2717 ? (n2366) : (n2710 ? (n2366) : (n2703 ? (n2366) : (n2696 ? (n2366) : (n2689 ? (n2366) : (n2682 ? (n2366) : (n2675 ? (n2366) : (n2668 ? (n2366) : (n2661 ? (n2366) : (n2654 ? (n2366) : (n2647 ? (n2366) : (n2640 ? (n2366) : (n2633 ? (n2366) : (n2626 ? (n2366) : (n2619 ? (n2366) : (n2612 ? (n2366) : (n2605 ? (n2366) : (n2598 ? (n2366) : (n2591 ? (n2366) : (n2584 ? (n2366) : (n2577 ? (n2366) : (n2570 ? (n2366) : (n2563 ? (n2366) : (n2556 ? (n2366) : (n2549 ? (n2366) : (n2542 ? (n2366) : (n2535 ? (n2366) : (n2528 ? (n2366) : (n2521 ? (n2366) : (n2514 ? (n2366) : (n2507 ? (n2366) : (n2500 ? (n2366) : (n2493 ? (n2366) : (n2486 ? (n2366) : (n2479 ? (n2366) : (n2472 ? (n2366) : (n2465 ? (n2366) : (n2458 ? (n2366) : (n2451 ? (n2366) : (n2444 ? (n2366) : (n2437 ? (n2366) : (n2430 ? (n2366) : (n2423 ? (n2366) : (n2416 ? (n2366) : (n2409 ? (n2366) : (n2402 ? (n2366) : (n2395 ? (n2366) : (n2388 ? (n2366) : (n2365 ? (n2366) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data0 = n3494 ? (n2367) : (n3487 ? (n2367) : (n3480 ? (n2367) : (n3473 ? (n2367) : (n3466 ? (n2367) : (n3459 ? (n2367) : (n3452 ? (n2367) : (n3445 ? (n2367) : (n3438 ? (n2367) : (n3431 ? (n2367) : (n3424 ? (n2367) : (n3417 ? (n2367) : (n3410 ? (n2367) : (n3403 ? (n2367) : (n3396 ? (n2367) : (n3389 ? (n2367) : (n3382 ? (n2367) : (n3375 ? (n2367) : (n3368 ? (n2367) : (n3361 ? (n2367) : (n3354 ? (n2367) : (n3347 ? (n2367) : (n3340 ? (n2367) : (n3333 ? (n2367) : (n3326 ? (n2367) : (n3319 ? (n2367) : (n3312 ? (n2367) : (n3305 ? (n2367) : (n3298 ? (n2367) : (n3291 ? (n2367) : (n3284 ? (n2367) : (n3277 ? (n2367) : (n3270 ? (n2367) : (n3263 ? (n2367) : (n3256 ? (n2367) : (n3249 ? (n2367) : (n3242 ? (n2367) : (n3235 ? (n2367) : (n3228 ? (n2367) : (n3221 ? (n2367) : (n3214 ? (n2367) : (n3207 ? (n2367) : (n3200 ? (n2367) : (n3193 ? (n2367) : (n3186 ? (n2367) : (n3179 ? (n2367) : (n3172 ? (n2367) : (n3165 ? (n2367) : (n3158 ? (n2367) : (n3151 ? (n2367) : (n3144 ? (n2367) : (n3137 ? (n2367) : (n3130 ? (n2367) : (n3123 ? (n2367) : (n3116 ? (n2367) : (n3109 ? (n2367) : (n3102 ? (n2367) : (n3095 ? (n2367) : (n3088 ? (n2367) : (n3081 ? (n2367) : (n3074 ? (n2367) : (n3067 ? (n2367) : (n3060 ? (n2367) : (n3053 ? (n2367) : (n3046 ? (n2367) : (n3039 ? (n2367) : (n3032 ? (n2367) : (n3025 ? (n2367) : (n3018 ? (n2367) : (n3011 ? (n2367) : (n3004 ? (n2367) : (n2997 ? (n2367) : (n2990 ? (n2367) : (n2983 ? (n2367) : (n2976 ? (n2367) : (n2969 ? (n2367) : (n2962 ? (n2367) : (n2955 ? (n2367) : (n2948 ? (n2367) : (n2941 ? (n2367) : (n2934 ? (n2367) : (n2927 ? (n2367) : (n2920 ? (n2367) : (n2913 ? (n2367) : (n2906 ? (n2367) : (n2899 ? (n2367) : (n2892 ? (n2367) : (n2885 ? (n2367) : (n2878 ? (n2367) : (n2871 ? (n2367) : (n2864 ? (n2367) : (n2857 ? (n2367) : (n2850 ? (n2367) : (n2843 ? (n2367) : (n2836 ? (n2367) : (n2829 ? (n2367) : (n2822 ? (n2367) : (n2815 ? (n2367) : (n2808 ? (n2367) : (n2801 ? (n2367) : (n2794 ? (n2367) : (n2787 ? (n2367) : (n2780 ? (n2367) : (n2773 ? (n2367) : (n2766 ? (n2367) : (n2759 ? (n2367) : (n2752 ? (n2367) : (n2745 ? (n2367) : (n2738 ? (n2367) : (n2731 ? (n2367) : (n2724 ? (n2367) : (n2717 ? (n2367) : (n2710 ? (n2367) : (n2703 ? (n2367) : (n2696 ? (n2367) : (n2689 ? (n2367) : (n2682 ? (n2367) : (n2675 ? (n2367) : (n2668 ? (n2367) : (n2661 ? (n2367) : (n2654 ? (n2367) : (n2647 ? (n2367) : (n2640 ? (n2367) : (n2633 ? (n2367) : (n2626 ? (n2367) : (n2619 ? (n2367) : (n2612 ? (n2367) : (n2605 ? (n2367) : (n2598 ? (n2367) : (n2591 ? (n2367) : (n2584 ? (n2367) : (n2577 ? (n2367) : (n2570 ? (n2367) : (n2563 ? (n2367) : (n2556 ? (n2367) : (n2549 ? (n2367) : (n2542 ? (n2367) : (n2535 ? (n2367) : (n2528 ? (n2367) : (n2521 ? (n2367) : (n2514 ? (n2367) : (n2507 ? (n2367) : (n2500 ? (n2367) : (n2493 ? (n2367) : (n2486 ? (n2367) : (n2479 ? (n2367) : (n2472 ? (n2367) : (n2465 ? (n2367) : (n2458 ? (n2367) : (n2451 ? (n2367) : (n2444 ? (n2367) : (n2437 ? (n2367) : (n2430 ? (n2367) : (n2423 ? (n2367) : (n2416 ? (n2367) : (n2409 ? (n2367) : (n2402 ? (n2367) : (n2395 ? (n2367) : (n2388 ? (n2367) : (n2365 ? (n2367) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen0 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr1 = n3494 ? (n2368) : (n3487 ? (n2368) : (n3480 ? (n2368) : (n3473 ? (n2368) : (n3466 ? (n2368) : (n3459 ? (n2368) : (n3452 ? (n2368) : (n3445 ? (n2368) : (n3438 ? (n2368) : (n3431 ? (n2368) : (n3424 ? (n2368) : (n3417 ? (n2368) : (n3410 ? (n2368) : (n3403 ? (n2368) : (n3396 ? (n2368) : (n3389 ? (n2368) : (n3382 ? (n2368) : (n3375 ? (n2368) : (n3368 ? (n2368) : (n3361 ? (n2368) : (n3354 ? (n2368) : (n3347 ? (n2368) : (n3340 ? (n2368) : (n3333 ? (n2368) : (n3326 ? (n2368) : (n3319 ? (n2368) : (n3312 ? (n2368) : (n3305 ? (n2368) : (n3298 ? (n2368) : (n3291 ? (n2368) : (n3284 ? (n2368) : (n3277 ? (n2368) : (n3270 ? (n2368) : (n3263 ? (n2368) : (n3256 ? (n2368) : (n3249 ? (n2368) : (n3242 ? (n2368) : (n3235 ? (n2368) : (n3228 ? (n2368) : (n3221 ? (n2368) : (n3214 ? (n2368) : (n3207 ? (n2368) : (n3200 ? (n2368) : (n3193 ? (n2368) : (n3186 ? (n2368) : (n3179 ? (n2368) : (n3172 ? (n2368) : (n3165 ? (n2368) : (n3158 ? (n2368) : (n3151 ? (n2368) : (n3144 ? (n2368) : (n3137 ? (n2368) : (n3130 ? (n2368) : (n3123 ? (n2368) : (n3116 ? (n2368) : (n3109 ? (n2368) : (n3102 ? (n2368) : (n3095 ? (n2368) : (n3088 ? (n2368) : (n3081 ? (n2368) : (n3074 ? (n2368) : (n3067 ? (n2368) : (n3060 ? (n2368) : (n3053 ? (n2368) : (n3046 ? (n2368) : (n3039 ? (n2368) : (n3032 ? (n2368) : (n3025 ? (n2368) : (n3018 ? (n2368) : (n3011 ? (n2368) : (n3004 ? (n2368) : (n2997 ? (n2368) : (n2990 ? (n2368) : (n2983 ? (n2368) : (n2976 ? (n2368) : (n2969 ? (n2368) : (n2962 ? (n2368) : (n2955 ? (n2368) : (n2948 ? (n2368) : (n2941 ? (n2368) : (n2934 ? (n2368) : (n2927 ? (n2368) : (n2920 ? (n2368) : (n2913 ? (n2368) : (n2906 ? (n2368) : (n2899 ? (n2368) : (n2892 ? (n2368) : (n2885 ? (n2368) : (n2878 ? (n2368) : (n2871 ? (n2368) : (n2864 ? (n2368) : (n2857 ? (n2368) : (n2850 ? (n2368) : (n2843 ? (n2368) : (n2836 ? (n2368) : (n2829 ? (n2368) : (n2822 ? (n2368) : (n2815 ? (n2368) : (n2808 ? (n2368) : (n2801 ? (n2368) : (n2794 ? (n2368) : (n2787 ? (n2368) : (n2780 ? (n2368) : (n2773 ? (n2368) : (n2766 ? (n2368) : (n2759 ? (n2368) : (n2752 ? (n2368) : (n2745 ? (n2368) : (n2738 ? (n2368) : (n2731 ? (n2368) : (n2724 ? (n2368) : (n2717 ? (n2368) : (n2710 ? (n2368) : (n2703 ? (n2368) : (n2696 ? (n2368) : (n2689 ? (n2368) : (n2682 ? (n2368) : (n2675 ? (n2368) : (n2668 ? (n2368) : (n2661 ? (n2368) : (n2654 ? (n2368) : (n2647 ? (n2368) : (n2640 ? (n2368) : (n2633 ? (n2368) : (n2626 ? (n2368) : (n2619 ? (n2368) : (n2612 ? (n2368) : (n2605 ? (n2368) : (n2598 ? (n2368) : (n2591 ? (n2368) : (n2584 ? (n2368) : (n2577 ? (n2368) : (n2570 ? (n2368) : (n2563 ? (n2368) : (n2556 ? (n2368) : (n2549 ? (n2368) : (n2542 ? (n2368) : (n2535 ? (n2368) : (n2528 ? (n2368) : (n2521 ? (n2368) : (n2514 ? (n2368) : (n2507 ? (n2368) : (n2500 ? (n2368) : (n2493 ? (n2368) : (n2486 ? (n2368) : (n2479 ? (n2368) : (n2472 ? (n2368) : (n2465 ? (n2368) : (n2458 ? (n2368) : (n2451 ? (n2368) : (n2444 ? (n2368) : (n2437 ? (n2368) : (n2430 ? (n2368) : (n2423 ? (n2368) : (n2416 ? (n2368) : (n2409 ? (n2368) : (n2402 ? (n2368) : (n2395 ? (n2368) : (n2388 ? (n2368) : (n2365 ? (n2368) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data1 = n3494 ? (n2369) : (n3487 ? (n2369) : (n3480 ? (n2369) : (n3473 ? (n2369) : (n3466 ? (n2369) : (n3459 ? (n2369) : (n3452 ? (n2369) : (n3445 ? (n2369) : (n3438 ? (n2369) : (n3431 ? (n2369) : (n3424 ? (n2369) : (n3417 ? (n2369) : (n3410 ? (n2369) : (n3403 ? (n2369) : (n3396 ? (n2369) : (n3389 ? (n2369) : (n3382 ? (n2369) : (n3375 ? (n2369) : (n3368 ? (n2369) : (n3361 ? (n2369) : (n3354 ? (n2369) : (n3347 ? (n2369) : (n3340 ? (n2369) : (n3333 ? (n2369) : (n3326 ? (n2369) : (n3319 ? (n2369) : (n3312 ? (n2369) : (n3305 ? (n2369) : (n3298 ? (n2369) : (n3291 ? (n2369) : (n3284 ? (n2369) : (n3277 ? (n2369) : (n3270 ? (n2369) : (n3263 ? (n2369) : (n3256 ? (n2369) : (n3249 ? (n2369) : (n3242 ? (n2369) : (n3235 ? (n2369) : (n3228 ? (n2369) : (n3221 ? (n2369) : (n3214 ? (n2369) : (n3207 ? (n2369) : (n3200 ? (n2369) : (n3193 ? (n2369) : (n3186 ? (n2369) : (n3179 ? (n2369) : (n3172 ? (n2369) : (n3165 ? (n2369) : (n3158 ? (n2369) : (n3151 ? (n2369) : (n3144 ? (n2369) : (n3137 ? (n2369) : (n3130 ? (n2369) : (n3123 ? (n2369) : (n3116 ? (n2369) : (n3109 ? (n2369) : (n3102 ? (n2369) : (n3095 ? (n2369) : (n3088 ? (n2369) : (n3081 ? (n2369) : (n3074 ? (n2369) : (n3067 ? (n2369) : (n3060 ? (n2369) : (n3053 ? (n2369) : (n3046 ? (n2369) : (n3039 ? (n2369) : (n3032 ? (n2369) : (n3025 ? (n2369) : (n3018 ? (n2369) : (n3011 ? (n2369) : (n3004 ? (n2369) : (n2997 ? (n2369) : (n2990 ? (n2369) : (n2983 ? (n2369) : (n2976 ? (n2369) : (n2969 ? (n2369) : (n2962 ? (n2369) : (n2955 ? (n2369) : (n2948 ? (n2369) : (n2941 ? (n2369) : (n2934 ? (n2369) : (n2927 ? (n2369) : (n2920 ? (n2369) : (n2913 ? (n2369) : (n2906 ? (n2369) : (n2899 ? (n2369) : (n2892 ? (n2369) : (n2885 ? (n2369) : (n2878 ? (n2369) : (n2871 ? (n2369) : (n2864 ? (n2369) : (n2857 ? (n2369) : (n2850 ? (n2369) : (n2843 ? (n2369) : (n2836 ? (n2369) : (n2829 ? (n2369) : (n2822 ? (n2369) : (n2815 ? (n2369) : (n2808 ? (n2369) : (n2801 ? (n2369) : (n2794 ? (n2369) : (n2787 ? (n2369) : (n2780 ? (n2369) : (n2773 ? (n2369) : (n2766 ? (n2369) : (n2759 ? (n2369) : (n2752 ? (n2369) : (n2745 ? (n2369) : (n2738 ? (n2369) : (n2731 ? (n2369) : (n2724 ? (n2369) : (n2717 ? (n2369) : (n2710 ? (n2369) : (n2703 ? (n2369) : (n2696 ? (n2369) : (n2689 ? (n2369) : (n2682 ? (n2369) : (n2675 ? (n2369) : (n2668 ? (n2369) : (n2661 ? (n2369) : (n2654 ? (n2369) : (n2647 ? (n2369) : (n2640 ? (n2369) : (n2633 ? (n2369) : (n2626 ? (n2369) : (n2619 ? (n2369) : (n2612 ? (n2369) : (n2605 ? (n2369) : (n2598 ? (n2369) : (n2591 ? (n2369) : (n2584 ? (n2369) : (n2577 ? (n2369) : (n2570 ? (n2369) : (n2563 ? (n2369) : (n2556 ? (n2369) : (n2549 ? (n2369) : (n2542 ? (n2369) : (n2535 ? (n2369) : (n2528 ? (n2369) : (n2521 ? (n2369) : (n2514 ? (n2369) : (n2507 ? (n2369) : (n2500 ? (n2369) : (n2493 ? (n2369) : (n2486 ? (n2369) : (n2479 ? (n2369) : (n2472 ? (n2369) : (n2465 ? (n2369) : (n2458 ? (n2369) : (n2451 ? (n2369) : (n2444 ? (n2369) : (n2437 ? (n2369) : (n2430 ? (n2369) : (n2423 ? (n2369) : (n2416 ? (n2369) : (n2409 ? (n2369) : (n2402 ? (n2369) : (n2395 ? (n2369) : (n2388 ? (n2369) : (n2365 ? (n2369) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen1 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr2 = n3494 ? (n2370) : (n3487 ? (n2370) : (n3480 ? (n2370) : (n3473 ? (n2370) : (n3466 ? (n2370) : (n3459 ? (n2370) : (n3452 ? (n2370) : (n3445 ? (n2370) : (n3438 ? (n2370) : (n3431 ? (n2370) : (n3424 ? (n2370) : (n3417 ? (n2370) : (n3410 ? (n2370) : (n3403 ? (n2370) : (n3396 ? (n2370) : (n3389 ? (n2370) : (n3382 ? (n2370) : (n3375 ? (n2370) : (n3368 ? (n2370) : (n3361 ? (n2370) : (n3354 ? (n2370) : (n3347 ? (n2370) : (n3340 ? (n2370) : (n3333 ? (n2370) : (n3326 ? (n2370) : (n3319 ? (n2370) : (n3312 ? (n2370) : (n3305 ? (n2370) : (n3298 ? (n2370) : (n3291 ? (n2370) : (n3284 ? (n2370) : (n3277 ? (n2370) : (n3270 ? (n2370) : (n3263 ? (n2370) : (n3256 ? (n2370) : (n3249 ? (n2370) : (n3242 ? (n2370) : (n3235 ? (n2370) : (n3228 ? (n2370) : (n3221 ? (n2370) : (n3214 ? (n2370) : (n3207 ? (n2370) : (n3200 ? (n2370) : (n3193 ? (n2370) : (n3186 ? (n2370) : (n3179 ? (n2370) : (n3172 ? (n2370) : (n3165 ? (n2370) : (n3158 ? (n2370) : (n3151 ? (n2370) : (n3144 ? (n2370) : (n3137 ? (n2370) : (n3130 ? (n2370) : (n3123 ? (n2370) : (n3116 ? (n2370) : (n3109 ? (n2370) : (n3102 ? (n2370) : (n3095 ? (n2370) : (n3088 ? (n2370) : (n3081 ? (n2370) : (n3074 ? (n2370) : (n3067 ? (n2370) : (n3060 ? (n2370) : (n3053 ? (n2370) : (n3046 ? (n2370) : (n3039 ? (n2370) : (n3032 ? (n2370) : (n3025 ? (n2370) : (n3018 ? (n2370) : (n3011 ? (n2370) : (n3004 ? (n2370) : (n2997 ? (n2370) : (n2990 ? (n2370) : (n2983 ? (n2370) : (n2976 ? (n2370) : (n2969 ? (n2370) : (n2962 ? (n2370) : (n2955 ? (n2370) : (n2948 ? (n2370) : (n2941 ? (n2370) : (n2934 ? (n2370) : (n2927 ? (n2370) : (n2920 ? (n2370) : (n2913 ? (n2370) : (n2906 ? (n2370) : (n2899 ? (n2370) : (n2892 ? (n2370) : (n2885 ? (n2370) : (n2878 ? (n2370) : (n2871 ? (n2370) : (n2864 ? (n2370) : (n2857 ? (n2370) : (n2850 ? (n2370) : (n2843 ? (n2370) : (n2836 ? (n2370) : (n2829 ? (n2370) : (n2822 ? (n2370) : (n2815 ? (n2370) : (n2808 ? (n2370) : (n2801 ? (n2370) : (n2794 ? (n2370) : (n2787 ? (n2370) : (n2780 ? (n2370) : (n2773 ? (n2370) : (n2766 ? (n2370) : (n2759 ? (n2370) : (n2752 ? (n2370) : (n2745 ? (n2370) : (n2738 ? (n2370) : (n2731 ? (n2370) : (n2724 ? (n2370) : (n2717 ? (n2370) : (n2710 ? (n2370) : (n2703 ? (n2370) : (n2696 ? (n2370) : (n2689 ? (n2370) : (n2682 ? (n2370) : (n2675 ? (n2370) : (n2668 ? (n2370) : (n2661 ? (n2370) : (n2654 ? (n2370) : (n2647 ? (n2370) : (n2640 ? (n2370) : (n2633 ? (n2370) : (n2626 ? (n2370) : (n2619 ? (n2370) : (n2612 ? (n2370) : (n2605 ? (n2370) : (n2598 ? (n2370) : (n2591 ? (n2370) : (n2584 ? (n2370) : (n2577 ? (n2370) : (n2570 ? (n2370) : (n2563 ? (n2370) : (n2556 ? (n2370) : (n2549 ? (n2370) : (n2542 ? (n2370) : (n2535 ? (n2370) : (n2528 ? (n2370) : (n2521 ? (n2370) : (n2514 ? (n2370) : (n2507 ? (n2370) : (n2500 ? (n2370) : (n2493 ? (n2370) : (n2486 ? (n2370) : (n2479 ? (n2370) : (n2472 ? (n2370) : (n2465 ? (n2370) : (n2458 ? (n2370) : (n2451 ? (n2370) : (n2444 ? (n2370) : (n2437 ? (n2370) : (n2430 ? (n2370) : (n2423 ? (n2370) : (n2416 ? (n2370) : (n2409 ? (n2370) : (n2402 ? (n2370) : (n2395 ? (n2370) : (n2388 ? (n2370) : (n2365 ? (n2370) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data2 = n3494 ? (n2371) : (n3487 ? (n2371) : (n3480 ? (n2371) : (n3473 ? (n2371) : (n3466 ? (n2371) : (n3459 ? (n2371) : (n3452 ? (n2371) : (n3445 ? (n2371) : (n3438 ? (n2371) : (n3431 ? (n2371) : (n3424 ? (n2371) : (n3417 ? (n2371) : (n3410 ? (n2371) : (n3403 ? (n2371) : (n3396 ? (n2371) : (n3389 ? (n2371) : (n3382 ? (n2371) : (n3375 ? (n2371) : (n3368 ? (n2371) : (n3361 ? (n2371) : (n3354 ? (n2371) : (n3347 ? (n2371) : (n3340 ? (n2371) : (n3333 ? (n2371) : (n3326 ? (n2371) : (n3319 ? (n2371) : (n3312 ? (n2371) : (n3305 ? (n2371) : (n3298 ? (n2371) : (n3291 ? (n2371) : (n3284 ? (n2371) : (n3277 ? (n2371) : (n3270 ? (n2371) : (n3263 ? (n2371) : (n3256 ? (n2371) : (n3249 ? (n2371) : (n3242 ? (n2371) : (n3235 ? (n2371) : (n3228 ? (n2371) : (n3221 ? (n2371) : (n3214 ? (n2371) : (n3207 ? (n2371) : (n3200 ? (n2371) : (n3193 ? (n2371) : (n3186 ? (n2371) : (n3179 ? (n2371) : (n3172 ? (n2371) : (n3165 ? (n2371) : (n3158 ? (n2371) : (n3151 ? (n2371) : (n3144 ? (n2371) : (n3137 ? (n2371) : (n3130 ? (n2371) : (n3123 ? (n2371) : (n3116 ? (n2371) : (n3109 ? (n2371) : (n3102 ? (n2371) : (n3095 ? (n2371) : (n3088 ? (n2371) : (n3081 ? (n2371) : (n3074 ? (n2371) : (n3067 ? (n2371) : (n3060 ? (n2371) : (n3053 ? (n2371) : (n3046 ? (n2371) : (n3039 ? (n2371) : (n3032 ? (n2371) : (n3025 ? (n2371) : (n3018 ? (n2371) : (n3011 ? (n2371) : (n3004 ? (n2371) : (n2997 ? (n2371) : (n2990 ? (n2371) : (n2983 ? (n2371) : (n2976 ? (n2371) : (n2969 ? (n2371) : (n2962 ? (n2371) : (n2955 ? (n2371) : (n2948 ? (n2371) : (n2941 ? (n2371) : (n2934 ? (n2371) : (n2927 ? (n2371) : (n2920 ? (n2371) : (n2913 ? (n2371) : (n2906 ? (n2371) : (n2899 ? (n2371) : (n2892 ? (n2371) : (n2885 ? (n2371) : (n2878 ? (n2371) : (n2871 ? (n2371) : (n2864 ? (n2371) : (n2857 ? (n2371) : (n2850 ? (n2371) : (n2843 ? (n2371) : (n2836 ? (n2371) : (n2829 ? (n2371) : (n2822 ? (n2371) : (n2815 ? (n2371) : (n2808 ? (n2371) : (n2801 ? (n2371) : (n2794 ? (n2371) : (n2787 ? (n2371) : (n2780 ? (n2371) : (n2773 ? (n2371) : (n2766 ? (n2371) : (n2759 ? (n2371) : (n2752 ? (n2371) : (n2745 ? (n2371) : (n2738 ? (n2371) : (n2731 ? (n2371) : (n2724 ? (n2371) : (n2717 ? (n2371) : (n2710 ? (n2371) : (n2703 ? (n2371) : (n2696 ? (n2371) : (n2689 ? (n2371) : (n2682 ? (n2371) : (n2675 ? (n2371) : (n2668 ? (n2371) : (n2661 ? (n2371) : (n2654 ? (n2371) : (n2647 ? (n2371) : (n2640 ? (n2371) : (n2633 ? (n2371) : (n2626 ? (n2371) : (n2619 ? (n2371) : (n2612 ? (n2371) : (n2605 ? (n2371) : (n2598 ? (n2371) : (n2591 ? (n2371) : (n2584 ? (n2371) : (n2577 ? (n2371) : (n2570 ? (n2371) : (n2563 ? (n2371) : (n2556 ? (n2371) : (n2549 ? (n2371) : (n2542 ? (n2371) : (n2535 ? (n2371) : (n2528 ? (n2371) : (n2521 ? (n2371) : (n2514 ? (n2371) : (n2507 ? (n2371) : (n2500 ? (n2371) : (n2493 ? (n2371) : (n2486 ? (n2371) : (n2479 ? (n2371) : (n2472 ? (n2371) : (n2465 ? (n2371) : (n2458 ? (n2371) : (n2451 ? (n2371) : (n2444 ? (n2371) : (n2437 ? (n2371) : (n2430 ? (n2371) : (n2423 ? (n2371) : (n2416 ? (n2371) : (n2409 ? (n2371) : (n2402 ? (n2371) : (n2395 ? (n2371) : (n2388 ? (n2371) : (n2365 ? (n2371) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen2 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr3 = n3494 ? (n2372) : (n3487 ? (n2372) : (n3480 ? (n2372) : (n3473 ? (n2372) : (n3466 ? (n2372) : (n3459 ? (n2372) : (n3452 ? (n2372) : (n3445 ? (n2372) : (n3438 ? (n2372) : (n3431 ? (n2372) : (n3424 ? (n2372) : (n3417 ? (n2372) : (n3410 ? (n2372) : (n3403 ? (n2372) : (n3396 ? (n2372) : (n3389 ? (n2372) : (n3382 ? (n2372) : (n3375 ? (n2372) : (n3368 ? (n2372) : (n3361 ? (n2372) : (n3354 ? (n2372) : (n3347 ? (n2372) : (n3340 ? (n2372) : (n3333 ? (n2372) : (n3326 ? (n2372) : (n3319 ? (n2372) : (n3312 ? (n2372) : (n3305 ? (n2372) : (n3298 ? (n2372) : (n3291 ? (n2372) : (n3284 ? (n2372) : (n3277 ? (n2372) : (n3270 ? (n2372) : (n3263 ? (n2372) : (n3256 ? (n2372) : (n3249 ? (n2372) : (n3242 ? (n2372) : (n3235 ? (n2372) : (n3228 ? (n2372) : (n3221 ? (n2372) : (n3214 ? (n2372) : (n3207 ? (n2372) : (n3200 ? (n2372) : (n3193 ? (n2372) : (n3186 ? (n2372) : (n3179 ? (n2372) : (n3172 ? (n2372) : (n3165 ? (n2372) : (n3158 ? (n2372) : (n3151 ? (n2372) : (n3144 ? (n2372) : (n3137 ? (n2372) : (n3130 ? (n2372) : (n3123 ? (n2372) : (n3116 ? (n2372) : (n3109 ? (n2372) : (n3102 ? (n2372) : (n3095 ? (n2372) : (n3088 ? (n2372) : (n3081 ? (n2372) : (n3074 ? (n2372) : (n3067 ? (n2372) : (n3060 ? (n2372) : (n3053 ? (n2372) : (n3046 ? (n2372) : (n3039 ? (n2372) : (n3032 ? (n2372) : (n3025 ? (n2372) : (n3018 ? (n2372) : (n3011 ? (n2372) : (n3004 ? (n2372) : (n2997 ? (n2372) : (n2990 ? (n2372) : (n2983 ? (n2372) : (n2976 ? (n2372) : (n2969 ? (n2372) : (n2962 ? (n2372) : (n2955 ? (n2372) : (n2948 ? (n2372) : (n2941 ? (n2372) : (n2934 ? (n2372) : (n2927 ? (n2372) : (n2920 ? (n2372) : (n2913 ? (n2372) : (n2906 ? (n2372) : (n2899 ? (n2372) : (n2892 ? (n2372) : (n2885 ? (n2372) : (n2878 ? (n2372) : (n2871 ? (n2372) : (n2864 ? (n2372) : (n2857 ? (n2372) : (n2850 ? (n2372) : (n2843 ? (n2372) : (n2836 ? (n2372) : (n2829 ? (n2372) : (n2822 ? (n2372) : (n2815 ? (n2372) : (n2808 ? (n2372) : (n2801 ? (n2372) : (n2794 ? (n2372) : (n2787 ? (n2372) : (n2780 ? (n2372) : (n2773 ? (n2372) : (n2766 ? (n2372) : (n2759 ? (n2372) : (n2752 ? (n2372) : (n2745 ? (n2372) : (n2738 ? (n2372) : (n2731 ? (n2372) : (n2724 ? (n2372) : (n2717 ? (n2372) : (n2710 ? (n2372) : (n2703 ? (n2372) : (n2696 ? (n2372) : (n2689 ? (n2372) : (n2682 ? (n2372) : (n2675 ? (n2372) : (n2668 ? (n2372) : (n2661 ? (n2372) : (n2654 ? (n2372) : (n2647 ? (n2372) : (n2640 ? (n2372) : (n2633 ? (n2372) : (n2626 ? (n2372) : (n2619 ? (n2372) : (n2612 ? (n2372) : (n2605 ? (n2372) : (n2598 ? (n2372) : (n2591 ? (n2372) : (n2584 ? (n2372) : (n2577 ? (n2372) : (n2570 ? (n2372) : (n2563 ? (n2372) : (n2556 ? (n2372) : (n2549 ? (n2372) : (n2542 ? (n2372) : (n2535 ? (n2372) : (n2528 ? (n2372) : (n2521 ? (n2372) : (n2514 ? (n2372) : (n2507 ? (n2372) : (n2500 ? (n2372) : (n2493 ? (n2372) : (n2486 ? (n2372) : (n2479 ? (n2372) : (n2472 ? (n2372) : (n2465 ? (n2372) : (n2458 ? (n2372) : (n2451 ? (n2372) : (n2444 ? (n2372) : (n2437 ? (n2372) : (n2430 ? (n2372) : (n2423 ? (n2372) : (n2416 ? (n2372) : (n2409 ? (n2372) : (n2402 ? (n2372) : (n2395 ? (n2372) : (n2388 ? (n2372) : (n2365 ? (n2372) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data3 = n3494 ? (n2373) : (n3487 ? (n2373) : (n3480 ? (n2373) : (n3473 ? (n2373) : (n3466 ? (n2373) : (n3459 ? (n2373) : (n3452 ? (n2373) : (n3445 ? (n2373) : (n3438 ? (n2373) : (n3431 ? (n2373) : (n3424 ? (n2373) : (n3417 ? (n2373) : (n3410 ? (n2373) : (n3403 ? (n2373) : (n3396 ? (n2373) : (n3389 ? (n2373) : (n3382 ? (n2373) : (n3375 ? (n2373) : (n3368 ? (n2373) : (n3361 ? (n2373) : (n3354 ? (n2373) : (n3347 ? (n2373) : (n3340 ? (n2373) : (n3333 ? (n2373) : (n3326 ? (n2373) : (n3319 ? (n2373) : (n3312 ? (n2373) : (n3305 ? (n2373) : (n3298 ? (n2373) : (n3291 ? (n2373) : (n3284 ? (n2373) : (n3277 ? (n2373) : (n3270 ? (n2373) : (n3263 ? (n2373) : (n3256 ? (n2373) : (n3249 ? (n2373) : (n3242 ? (n2373) : (n3235 ? (n2373) : (n3228 ? (n2373) : (n3221 ? (n2373) : (n3214 ? (n2373) : (n3207 ? (n2373) : (n3200 ? (n2373) : (n3193 ? (n2373) : (n3186 ? (n2373) : (n3179 ? (n2373) : (n3172 ? (n2373) : (n3165 ? (n2373) : (n3158 ? (n2373) : (n3151 ? (n2373) : (n3144 ? (n2373) : (n3137 ? (n2373) : (n3130 ? (n2373) : (n3123 ? (n2373) : (n3116 ? (n2373) : (n3109 ? (n2373) : (n3102 ? (n2373) : (n3095 ? (n2373) : (n3088 ? (n2373) : (n3081 ? (n2373) : (n3074 ? (n2373) : (n3067 ? (n2373) : (n3060 ? (n2373) : (n3053 ? (n2373) : (n3046 ? (n2373) : (n3039 ? (n2373) : (n3032 ? (n2373) : (n3025 ? (n2373) : (n3018 ? (n2373) : (n3011 ? (n2373) : (n3004 ? (n2373) : (n2997 ? (n2373) : (n2990 ? (n2373) : (n2983 ? (n2373) : (n2976 ? (n2373) : (n2969 ? (n2373) : (n2962 ? (n2373) : (n2955 ? (n2373) : (n2948 ? (n2373) : (n2941 ? (n2373) : (n2934 ? (n2373) : (n2927 ? (n2373) : (n2920 ? (n2373) : (n2913 ? (n2373) : (n2906 ? (n2373) : (n2899 ? (n2373) : (n2892 ? (n2373) : (n2885 ? (n2373) : (n2878 ? (n2373) : (n2871 ? (n2373) : (n2864 ? (n2373) : (n2857 ? (n2373) : (n2850 ? (n2373) : (n2843 ? (n2373) : (n2836 ? (n2373) : (n2829 ? (n2373) : (n2822 ? (n2373) : (n2815 ? (n2373) : (n2808 ? (n2373) : (n2801 ? (n2373) : (n2794 ? (n2373) : (n2787 ? (n2373) : (n2780 ? (n2373) : (n2773 ? (n2373) : (n2766 ? (n2373) : (n2759 ? (n2373) : (n2752 ? (n2373) : (n2745 ? (n2373) : (n2738 ? (n2373) : (n2731 ? (n2373) : (n2724 ? (n2373) : (n2717 ? (n2373) : (n2710 ? (n2373) : (n2703 ? (n2373) : (n2696 ? (n2373) : (n2689 ? (n2373) : (n2682 ? (n2373) : (n2675 ? (n2373) : (n2668 ? (n2373) : (n2661 ? (n2373) : (n2654 ? (n2373) : (n2647 ? (n2373) : (n2640 ? (n2373) : (n2633 ? (n2373) : (n2626 ? (n2373) : (n2619 ? (n2373) : (n2612 ? (n2373) : (n2605 ? (n2373) : (n2598 ? (n2373) : (n2591 ? (n2373) : (n2584 ? (n2373) : (n2577 ? (n2373) : (n2570 ? (n2373) : (n2563 ? (n2373) : (n2556 ? (n2373) : (n2549 ? (n2373) : (n2542 ? (n2373) : (n2535 ? (n2373) : (n2528 ? (n2373) : (n2521 ? (n2373) : (n2514 ? (n2373) : (n2507 ? (n2373) : (n2500 ? (n2373) : (n2493 ? (n2373) : (n2486 ? (n2373) : (n2479 ? (n2373) : (n2472 ? (n2373) : (n2465 ? (n2373) : (n2458 ? (n2373) : (n2451 ? (n2373) : (n2444 ? (n2373) : (n2437 ? (n2373) : (n2430 ? (n2373) : (n2423 ? (n2373) : (n2416 ? (n2373) : (n2409 ? (n2373) : (n2402 ? (n2373) : (n2395 ? (n2373) : (n2388 ? (n2373) : (n2365 ? (n2373) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen3 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr4 = n3494 ? (n2374) : (n3487 ? (n2374) : (n3480 ? (n2374) : (n3473 ? (n2374) : (n3466 ? (n2374) : (n3459 ? (n2374) : (n3452 ? (n2374) : (n3445 ? (n2374) : (n3438 ? (n2374) : (n3431 ? (n2374) : (n3424 ? (n2374) : (n3417 ? (n2374) : (n3410 ? (n2374) : (n3403 ? (n2374) : (n3396 ? (n2374) : (n3389 ? (n2374) : (n3382 ? (n2374) : (n3375 ? (n2374) : (n3368 ? (n2374) : (n3361 ? (n2374) : (n3354 ? (n2374) : (n3347 ? (n2374) : (n3340 ? (n2374) : (n3333 ? (n2374) : (n3326 ? (n2374) : (n3319 ? (n2374) : (n3312 ? (n2374) : (n3305 ? (n2374) : (n3298 ? (n2374) : (n3291 ? (n2374) : (n3284 ? (n2374) : (n3277 ? (n2374) : (n3270 ? (n2374) : (n3263 ? (n2374) : (n3256 ? (n2374) : (n3249 ? (n2374) : (n3242 ? (n2374) : (n3235 ? (n2374) : (n3228 ? (n2374) : (n3221 ? (n2374) : (n3214 ? (n2374) : (n3207 ? (n2374) : (n3200 ? (n2374) : (n3193 ? (n2374) : (n3186 ? (n2374) : (n3179 ? (n2374) : (n3172 ? (n2374) : (n3165 ? (n2374) : (n3158 ? (n2374) : (n3151 ? (n2374) : (n3144 ? (n2374) : (n3137 ? (n2374) : (n3130 ? (n2374) : (n3123 ? (n2374) : (n3116 ? (n2374) : (n3109 ? (n2374) : (n3102 ? (n2374) : (n3095 ? (n2374) : (n3088 ? (n2374) : (n3081 ? (n2374) : (n3074 ? (n2374) : (n3067 ? (n2374) : (n3060 ? (n2374) : (n3053 ? (n2374) : (n3046 ? (n2374) : (n3039 ? (n2374) : (n3032 ? (n2374) : (n3025 ? (n2374) : (n3018 ? (n2374) : (n3011 ? (n2374) : (n3004 ? (n2374) : (n2997 ? (n2374) : (n2990 ? (n2374) : (n2983 ? (n2374) : (n2976 ? (n2374) : (n2969 ? (n2374) : (n2962 ? (n2374) : (n2955 ? (n2374) : (n2948 ? (n2374) : (n2941 ? (n2374) : (n2934 ? (n2374) : (n2927 ? (n2374) : (n2920 ? (n2374) : (n2913 ? (n2374) : (n2906 ? (n2374) : (n2899 ? (n2374) : (n2892 ? (n2374) : (n2885 ? (n2374) : (n2878 ? (n2374) : (n2871 ? (n2374) : (n2864 ? (n2374) : (n2857 ? (n2374) : (n2850 ? (n2374) : (n2843 ? (n2374) : (n2836 ? (n2374) : (n2829 ? (n2374) : (n2822 ? (n2374) : (n2815 ? (n2374) : (n2808 ? (n2374) : (n2801 ? (n2374) : (n2794 ? (n2374) : (n2787 ? (n2374) : (n2780 ? (n2374) : (n2773 ? (n2374) : (n2766 ? (n2374) : (n2759 ? (n2374) : (n2752 ? (n2374) : (n2745 ? (n2374) : (n2738 ? (n2374) : (n2731 ? (n2374) : (n2724 ? (n2374) : (n2717 ? (n2374) : (n2710 ? (n2374) : (n2703 ? (n2374) : (n2696 ? (n2374) : (n2689 ? (n2374) : (n2682 ? (n2374) : (n2675 ? (n2374) : (n2668 ? (n2374) : (n2661 ? (n2374) : (n2654 ? (n2374) : (n2647 ? (n2374) : (n2640 ? (n2374) : (n2633 ? (n2374) : (n2626 ? (n2374) : (n2619 ? (n2374) : (n2612 ? (n2374) : (n2605 ? (n2374) : (n2598 ? (n2374) : (n2591 ? (n2374) : (n2584 ? (n2374) : (n2577 ? (n2374) : (n2570 ? (n2374) : (n2563 ? (n2374) : (n2556 ? (n2374) : (n2549 ? (n2374) : (n2542 ? (n2374) : (n2535 ? (n2374) : (n2528 ? (n2374) : (n2521 ? (n2374) : (n2514 ? (n2374) : (n2507 ? (n2374) : (n2500 ? (n2374) : (n2493 ? (n2374) : (n2486 ? (n2374) : (n2479 ? (n2374) : (n2472 ? (n2374) : (n2465 ? (n2374) : (n2458 ? (n2374) : (n2451 ? (n2374) : (n2444 ? (n2374) : (n2437 ? (n2374) : (n2430 ? (n2374) : (n2423 ? (n2374) : (n2416 ? (n2374) : (n2409 ? (n2374) : (n2402 ? (n2374) : (n2395 ? (n2374) : (n2388 ? (n2374) : (n2365 ? (n2374) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data4 = n3494 ? (n2375) : (n3487 ? (n2375) : (n3480 ? (n2375) : (n3473 ? (n2375) : (n3466 ? (n2375) : (n3459 ? (n2375) : (n3452 ? (n2375) : (n3445 ? (n2375) : (n3438 ? (n2375) : (n3431 ? (n2375) : (n3424 ? (n2375) : (n3417 ? (n2375) : (n3410 ? (n2375) : (n3403 ? (n2375) : (n3396 ? (n2375) : (n3389 ? (n2375) : (n3382 ? (n2375) : (n3375 ? (n2375) : (n3368 ? (n2375) : (n3361 ? (n2375) : (n3354 ? (n2375) : (n3347 ? (n2375) : (n3340 ? (n2375) : (n3333 ? (n2375) : (n3326 ? (n2375) : (n3319 ? (n2375) : (n3312 ? (n2375) : (n3305 ? (n2375) : (n3298 ? (n2375) : (n3291 ? (n2375) : (n3284 ? (n2375) : (n3277 ? (n2375) : (n3270 ? (n2375) : (n3263 ? (n2375) : (n3256 ? (n2375) : (n3249 ? (n2375) : (n3242 ? (n2375) : (n3235 ? (n2375) : (n3228 ? (n2375) : (n3221 ? (n2375) : (n3214 ? (n2375) : (n3207 ? (n2375) : (n3200 ? (n2375) : (n3193 ? (n2375) : (n3186 ? (n2375) : (n3179 ? (n2375) : (n3172 ? (n2375) : (n3165 ? (n2375) : (n3158 ? (n2375) : (n3151 ? (n2375) : (n3144 ? (n2375) : (n3137 ? (n2375) : (n3130 ? (n2375) : (n3123 ? (n2375) : (n3116 ? (n2375) : (n3109 ? (n2375) : (n3102 ? (n2375) : (n3095 ? (n2375) : (n3088 ? (n2375) : (n3081 ? (n2375) : (n3074 ? (n2375) : (n3067 ? (n2375) : (n3060 ? (n2375) : (n3053 ? (n2375) : (n3046 ? (n2375) : (n3039 ? (n2375) : (n3032 ? (n2375) : (n3025 ? (n2375) : (n3018 ? (n2375) : (n3011 ? (n2375) : (n3004 ? (n2375) : (n2997 ? (n2375) : (n2990 ? (n2375) : (n2983 ? (n2375) : (n2976 ? (n2375) : (n2969 ? (n2375) : (n2962 ? (n2375) : (n2955 ? (n2375) : (n2948 ? (n2375) : (n2941 ? (n2375) : (n2934 ? (n2375) : (n2927 ? (n2375) : (n2920 ? (n2375) : (n2913 ? (n2375) : (n2906 ? (n2375) : (n2899 ? (n2375) : (n2892 ? (n2375) : (n2885 ? (n2375) : (n2878 ? (n2375) : (n2871 ? (n2375) : (n2864 ? (n2375) : (n2857 ? (n2375) : (n2850 ? (n2375) : (n2843 ? (n2375) : (n2836 ? (n2375) : (n2829 ? (n2375) : (n2822 ? (n2375) : (n2815 ? (n2375) : (n2808 ? (n2375) : (n2801 ? (n2375) : (n2794 ? (n2375) : (n2787 ? (n2375) : (n2780 ? (n2375) : (n2773 ? (n2375) : (n2766 ? (n2375) : (n2759 ? (n2375) : (n2752 ? (n2375) : (n2745 ? (n2375) : (n2738 ? (n2375) : (n2731 ? (n2375) : (n2724 ? (n2375) : (n2717 ? (n2375) : (n2710 ? (n2375) : (n2703 ? (n2375) : (n2696 ? (n2375) : (n2689 ? (n2375) : (n2682 ? (n2375) : (n2675 ? (n2375) : (n2668 ? (n2375) : (n2661 ? (n2375) : (n2654 ? (n2375) : (n2647 ? (n2375) : (n2640 ? (n2375) : (n2633 ? (n2375) : (n2626 ? (n2375) : (n2619 ? (n2375) : (n2612 ? (n2375) : (n2605 ? (n2375) : (n2598 ? (n2375) : (n2591 ? (n2375) : (n2584 ? (n2375) : (n2577 ? (n2375) : (n2570 ? (n2375) : (n2563 ? (n2375) : (n2556 ? (n2375) : (n2549 ? (n2375) : (n2542 ? (n2375) : (n2535 ? (n2375) : (n2528 ? (n2375) : (n2521 ? (n2375) : (n2514 ? (n2375) : (n2507 ? (n2375) : (n2500 ? (n2375) : (n2493 ? (n2375) : (n2486 ? (n2375) : (n2479 ? (n2375) : (n2472 ? (n2375) : (n2465 ? (n2375) : (n2458 ? (n2375) : (n2451 ? (n2375) : (n2444 ? (n2375) : (n2437 ? (n2375) : (n2430 ? (n2375) : (n2423 ? (n2375) : (n2416 ? (n2375) : (n2409 ? (n2375) : (n2402 ? (n2375) : (n2395 ? (n2375) : (n2388 ? (n2375) : (n2365 ? (n2375) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen4 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr5 = n3494 ? (n2376) : (n3487 ? (n2376) : (n3480 ? (n2376) : (n3473 ? (n2376) : (n3466 ? (n2376) : (n3459 ? (n2376) : (n3452 ? (n2376) : (n3445 ? (n2376) : (n3438 ? (n2376) : (n3431 ? (n2376) : (n3424 ? (n2376) : (n3417 ? (n2376) : (n3410 ? (n2376) : (n3403 ? (n2376) : (n3396 ? (n2376) : (n3389 ? (n2376) : (n3382 ? (n2376) : (n3375 ? (n2376) : (n3368 ? (n2376) : (n3361 ? (n2376) : (n3354 ? (n2376) : (n3347 ? (n2376) : (n3340 ? (n2376) : (n3333 ? (n2376) : (n3326 ? (n2376) : (n3319 ? (n2376) : (n3312 ? (n2376) : (n3305 ? (n2376) : (n3298 ? (n2376) : (n3291 ? (n2376) : (n3284 ? (n2376) : (n3277 ? (n2376) : (n3270 ? (n2376) : (n3263 ? (n2376) : (n3256 ? (n2376) : (n3249 ? (n2376) : (n3242 ? (n2376) : (n3235 ? (n2376) : (n3228 ? (n2376) : (n3221 ? (n2376) : (n3214 ? (n2376) : (n3207 ? (n2376) : (n3200 ? (n2376) : (n3193 ? (n2376) : (n3186 ? (n2376) : (n3179 ? (n2376) : (n3172 ? (n2376) : (n3165 ? (n2376) : (n3158 ? (n2376) : (n3151 ? (n2376) : (n3144 ? (n2376) : (n3137 ? (n2376) : (n3130 ? (n2376) : (n3123 ? (n2376) : (n3116 ? (n2376) : (n3109 ? (n2376) : (n3102 ? (n2376) : (n3095 ? (n2376) : (n3088 ? (n2376) : (n3081 ? (n2376) : (n3074 ? (n2376) : (n3067 ? (n2376) : (n3060 ? (n2376) : (n3053 ? (n2376) : (n3046 ? (n2376) : (n3039 ? (n2376) : (n3032 ? (n2376) : (n3025 ? (n2376) : (n3018 ? (n2376) : (n3011 ? (n2376) : (n3004 ? (n2376) : (n2997 ? (n2376) : (n2990 ? (n2376) : (n2983 ? (n2376) : (n2976 ? (n2376) : (n2969 ? (n2376) : (n2962 ? (n2376) : (n2955 ? (n2376) : (n2948 ? (n2376) : (n2941 ? (n2376) : (n2934 ? (n2376) : (n2927 ? (n2376) : (n2920 ? (n2376) : (n2913 ? (n2376) : (n2906 ? (n2376) : (n2899 ? (n2376) : (n2892 ? (n2376) : (n2885 ? (n2376) : (n2878 ? (n2376) : (n2871 ? (n2376) : (n2864 ? (n2376) : (n2857 ? (n2376) : (n2850 ? (n2376) : (n2843 ? (n2376) : (n2836 ? (n2376) : (n2829 ? (n2376) : (n2822 ? (n2376) : (n2815 ? (n2376) : (n2808 ? (n2376) : (n2801 ? (n2376) : (n2794 ? (n2376) : (n2787 ? (n2376) : (n2780 ? (n2376) : (n2773 ? (n2376) : (n2766 ? (n2376) : (n2759 ? (n2376) : (n2752 ? (n2376) : (n2745 ? (n2376) : (n2738 ? (n2376) : (n2731 ? (n2376) : (n2724 ? (n2376) : (n2717 ? (n2376) : (n2710 ? (n2376) : (n2703 ? (n2376) : (n2696 ? (n2376) : (n2689 ? (n2376) : (n2682 ? (n2376) : (n2675 ? (n2376) : (n2668 ? (n2376) : (n2661 ? (n2376) : (n2654 ? (n2376) : (n2647 ? (n2376) : (n2640 ? (n2376) : (n2633 ? (n2376) : (n2626 ? (n2376) : (n2619 ? (n2376) : (n2612 ? (n2376) : (n2605 ? (n2376) : (n2598 ? (n2376) : (n2591 ? (n2376) : (n2584 ? (n2376) : (n2577 ? (n2376) : (n2570 ? (n2376) : (n2563 ? (n2376) : (n2556 ? (n2376) : (n2549 ? (n2376) : (n2542 ? (n2376) : (n2535 ? (n2376) : (n2528 ? (n2376) : (n2521 ? (n2376) : (n2514 ? (n2376) : (n2507 ? (n2376) : (n2500 ? (n2376) : (n2493 ? (n2376) : (n2486 ? (n2376) : (n2479 ? (n2376) : (n2472 ? (n2376) : (n2465 ? (n2376) : (n2458 ? (n2376) : (n2451 ? (n2376) : (n2444 ? (n2376) : (n2437 ? (n2376) : (n2430 ? (n2376) : (n2423 ? (n2376) : (n2416 ? (n2376) : (n2409 ? (n2376) : (n2402 ? (n2376) : (n2395 ? (n2376) : (n2388 ? (n2376) : (n2365 ? (n2376) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data5 = n3494 ? (n2377) : (n3487 ? (n2377) : (n3480 ? (n2377) : (n3473 ? (n2377) : (n3466 ? (n2377) : (n3459 ? (n2377) : (n3452 ? (n2377) : (n3445 ? (n2377) : (n3438 ? (n2377) : (n3431 ? (n2377) : (n3424 ? (n2377) : (n3417 ? (n2377) : (n3410 ? (n2377) : (n3403 ? (n2377) : (n3396 ? (n2377) : (n3389 ? (n2377) : (n3382 ? (n2377) : (n3375 ? (n2377) : (n3368 ? (n2377) : (n3361 ? (n2377) : (n3354 ? (n2377) : (n3347 ? (n2377) : (n3340 ? (n2377) : (n3333 ? (n2377) : (n3326 ? (n2377) : (n3319 ? (n2377) : (n3312 ? (n2377) : (n3305 ? (n2377) : (n3298 ? (n2377) : (n3291 ? (n2377) : (n3284 ? (n2377) : (n3277 ? (n2377) : (n3270 ? (n2377) : (n3263 ? (n2377) : (n3256 ? (n2377) : (n3249 ? (n2377) : (n3242 ? (n2377) : (n3235 ? (n2377) : (n3228 ? (n2377) : (n3221 ? (n2377) : (n3214 ? (n2377) : (n3207 ? (n2377) : (n3200 ? (n2377) : (n3193 ? (n2377) : (n3186 ? (n2377) : (n3179 ? (n2377) : (n3172 ? (n2377) : (n3165 ? (n2377) : (n3158 ? (n2377) : (n3151 ? (n2377) : (n3144 ? (n2377) : (n3137 ? (n2377) : (n3130 ? (n2377) : (n3123 ? (n2377) : (n3116 ? (n2377) : (n3109 ? (n2377) : (n3102 ? (n2377) : (n3095 ? (n2377) : (n3088 ? (n2377) : (n3081 ? (n2377) : (n3074 ? (n2377) : (n3067 ? (n2377) : (n3060 ? (n2377) : (n3053 ? (n2377) : (n3046 ? (n2377) : (n3039 ? (n2377) : (n3032 ? (n2377) : (n3025 ? (n2377) : (n3018 ? (n2377) : (n3011 ? (n2377) : (n3004 ? (n2377) : (n2997 ? (n2377) : (n2990 ? (n2377) : (n2983 ? (n2377) : (n2976 ? (n2377) : (n2969 ? (n2377) : (n2962 ? (n2377) : (n2955 ? (n2377) : (n2948 ? (n2377) : (n2941 ? (n2377) : (n2934 ? (n2377) : (n2927 ? (n2377) : (n2920 ? (n2377) : (n2913 ? (n2377) : (n2906 ? (n2377) : (n2899 ? (n2377) : (n2892 ? (n2377) : (n2885 ? (n2377) : (n2878 ? (n2377) : (n2871 ? (n2377) : (n2864 ? (n2377) : (n2857 ? (n2377) : (n2850 ? (n2377) : (n2843 ? (n2377) : (n2836 ? (n2377) : (n2829 ? (n2377) : (n2822 ? (n2377) : (n2815 ? (n2377) : (n2808 ? (n2377) : (n2801 ? (n2377) : (n2794 ? (n2377) : (n2787 ? (n2377) : (n2780 ? (n2377) : (n2773 ? (n2377) : (n2766 ? (n2377) : (n2759 ? (n2377) : (n2752 ? (n2377) : (n2745 ? (n2377) : (n2738 ? (n2377) : (n2731 ? (n2377) : (n2724 ? (n2377) : (n2717 ? (n2377) : (n2710 ? (n2377) : (n2703 ? (n2377) : (n2696 ? (n2377) : (n2689 ? (n2377) : (n2682 ? (n2377) : (n2675 ? (n2377) : (n2668 ? (n2377) : (n2661 ? (n2377) : (n2654 ? (n2377) : (n2647 ? (n2377) : (n2640 ? (n2377) : (n2633 ? (n2377) : (n2626 ? (n2377) : (n2619 ? (n2377) : (n2612 ? (n2377) : (n2605 ? (n2377) : (n2598 ? (n2377) : (n2591 ? (n2377) : (n2584 ? (n2377) : (n2577 ? (n2377) : (n2570 ? (n2377) : (n2563 ? (n2377) : (n2556 ? (n2377) : (n2549 ? (n2377) : (n2542 ? (n2377) : (n2535 ? (n2377) : (n2528 ? (n2377) : (n2521 ? (n2377) : (n2514 ? (n2377) : (n2507 ? (n2377) : (n2500 ? (n2377) : (n2493 ? (n2377) : (n2486 ? (n2377) : (n2479 ? (n2377) : (n2472 ? (n2377) : (n2465 ? (n2377) : (n2458 ? (n2377) : (n2451 ? (n2377) : (n2444 ? (n2377) : (n2437 ? (n2377) : (n2430 ? (n2377) : (n2423 ? (n2377) : (n2416 ? (n2377) : (n2409 ? (n2377) : (n2402 ? (n2377) : (n2395 ? (n2377) : (n2388 ? (n2377) : (n2365 ? (n2377) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen5 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr6 = n3494 ? (n2378) : (n3487 ? (n2378) : (n3480 ? (n2378) : (n3473 ? (n2378) : (n3466 ? (n2378) : (n3459 ? (n2378) : (n3452 ? (n2378) : (n3445 ? (n2378) : (n3438 ? (n2378) : (n3431 ? (n2378) : (n3424 ? (n2378) : (n3417 ? (n2378) : (n3410 ? (n2378) : (n3403 ? (n2378) : (n3396 ? (n2378) : (n3389 ? (n2378) : (n3382 ? (n2378) : (n3375 ? (n2378) : (n3368 ? (n2378) : (n3361 ? (n2378) : (n3354 ? (n2378) : (n3347 ? (n2378) : (n3340 ? (n2378) : (n3333 ? (n2378) : (n3326 ? (n2378) : (n3319 ? (n2378) : (n3312 ? (n2378) : (n3305 ? (n2378) : (n3298 ? (n2378) : (n3291 ? (n2378) : (n3284 ? (n2378) : (n3277 ? (n2378) : (n3270 ? (n2378) : (n3263 ? (n2378) : (n3256 ? (n2378) : (n3249 ? (n2378) : (n3242 ? (n2378) : (n3235 ? (n2378) : (n3228 ? (n2378) : (n3221 ? (n2378) : (n3214 ? (n2378) : (n3207 ? (n2378) : (n3200 ? (n2378) : (n3193 ? (n2378) : (n3186 ? (n2378) : (n3179 ? (n2378) : (n3172 ? (n2378) : (n3165 ? (n2378) : (n3158 ? (n2378) : (n3151 ? (n2378) : (n3144 ? (n2378) : (n3137 ? (n2378) : (n3130 ? (n2378) : (n3123 ? (n2378) : (n3116 ? (n2378) : (n3109 ? (n2378) : (n3102 ? (n2378) : (n3095 ? (n2378) : (n3088 ? (n2378) : (n3081 ? (n2378) : (n3074 ? (n2378) : (n3067 ? (n2378) : (n3060 ? (n2378) : (n3053 ? (n2378) : (n3046 ? (n2378) : (n3039 ? (n2378) : (n3032 ? (n2378) : (n3025 ? (n2378) : (n3018 ? (n2378) : (n3011 ? (n2378) : (n3004 ? (n2378) : (n2997 ? (n2378) : (n2990 ? (n2378) : (n2983 ? (n2378) : (n2976 ? (n2378) : (n2969 ? (n2378) : (n2962 ? (n2378) : (n2955 ? (n2378) : (n2948 ? (n2378) : (n2941 ? (n2378) : (n2934 ? (n2378) : (n2927 ? (n2378) : (n2920 ? (n2378) : (n2913 ? (n2378) : (n2906 ? (n2378) : (n2899 ? (n2378) : (n2892 ? (n2378) : (n2885 ? (n2378) : (n2878 ? (n2378) : (n2871 ? (n2378) : (n2864 ? (n2378) : (n2857 ? (n2378) : (n2850 ? (n2378) : (n2843 ? (n2378) : (n2836 ? (n2378) : (n2829 ? (n2378) : (n2822 ? (n2378) : (n2815 ? (n2378) : (n2808 ? (n2378) : (n2801 ? (n2378) : (n2794 ? (n2378) : (n2787 ? (n2378) : (n2780 ? (n2378) : (n2773 ? (n2378) : (n2766 ? (n2378) : (n2759 ? (n2378) : (n2752 ? (n2378) : (n2745 ? (n2378) : (n2738 ? (n2378) : (n2731 ? (n2378) : (n2724 ? (n2378) : (n2717 ? (n2378) : (n2710 ? (n2378) : (n2703 ? (n2378) : (n2696 ? (n2378) : (n2689 ? (n2378) : (n2682 ? (n2378) : (n2675 ? (n2378) : (n2668 ? (n2378) : (n2661 ? (n2378) : (n2654 ? (n2378) : (n2647 ? (n2378) : (n2640 ? (n2378) : (n2633 ? (n2378) : (n2626 ? (n2378) : (n2619 ? (n2378) : (n2612 ? (n2378) : (n2605 ? (n2378) : (n2598 ? (n2378) : (n2591 ? (n2378) : (n2584 ? (n2378) : (n2577 ? (n2378) : (n2570 ? (n2378) : (n2563 ? (n2378) : (n2556 ? (n2378) : (n2549 ? (n2378) : (n2542 ? (n2378) : (n2535 ? (n2378) : (n2528 ? (n2378) : (n2521 ? (n2378) : (n2514 ? (n2378) : (n2507 ? (n2378) : (n2500 ? (n2378) : (n2493 ? (n2378) : (n2486 ? (n2378) : (n2479 ? (n2378) : (n2472 ? (n2378) : (n2465 ? (n2378) : (n2458 ? (n2378) : (n2451 ? (n2378) : (n2444 ? (n2378) : (n2437 ? (n2378) : (n2430 ? (n2378) : (n2423 ? (n2378) : (n2416 ? (n2378) : (n2409 ? (n2378) : (n2402 ? (n2378) : (n2395 ? (n2378) : (n2388 ? (n2378) : (n2365 ? (n2378) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data6 = n3494 ? (n2379) : (n3487 ? (n2379) : (n3480 ? (n2379) : (n3473 ? (n2379) : (n3466 ? (n2379) : (n3459 ? (n2379) : (n3452 ? (n2379) : (n3445 ? (n2379) : (n3438 ? (n2379) : (n3431 ? (n2379) : (n3424 ? (n2379) : (n3417 ? (n2379) : (n3410 ? (n2379) : (n3403 ? (n2379) : (n3396 ? (n2379) : (n3389 ? (n2379) : (n3382 ? (n2379) : (n3375 ? (n2379) : (n3368 ? (n2379) : (n3361 ? (n2379) : (n3354 ? (n2379) : (n3347 ? (n2379) : (n3340 ? (n2379) : (n3333 ? (n2379) : (n3326 ? (n2379) : (n3319 ? (n2379) : (n3312 ? (n2379) : (n3305 ? (n2379) : (n3298 ? (n2379) : (n3291 ? (n2379) : (n3284 ? (n2379) : (n3277 ? (n2379) : (n3270 ? (n2379) : (n3263 ? (n2379) : (n3256 ? (n2379) : (n3249 ? (n2379) : (n3242 ? (n2379) : (n3235 ? (n2379) : (n3228 ? (n2379) : (n3221 ? (n2379) : (n3214 ? (n2379) : (n3207 ? (n2379) : (n3200 ? (n2379) : (n3193 ? (n2379) : (n3186 ? (n2379) : (n3179 ? (n2379) : (n3172 ? (n2379) : (n3165 ? (n2379) : (n3158 ? (n2379) : (n3151 ? (n2379) : (n3144 ? (n2379) : (n3137 ? (n2379) : (n3130 ? (n2379) : (n3123 ? (n2379) : (n3116 ? (n2379) : (n3109 ? (n2379) : (n3102 ? (n2379) : (n3095 ? (n2379) : (n3088 ? (n2379) : (n3081 ? (n2379) : (n3074 ? (n2379) : (n3067 ? (n2379) : (n3060 ? (n2379) : (n3053 ? (n2379) : (n3046 ? (n2379) : (n3039 ? (n2379) : (n3032 ? (n2379) : (n3025 ? (n2379) : (n3018 ? (n2379) : (n3011 ? (n2379) : (n3004 ? (n2379) : (n2997 ? (n2379) : (n2990 ? (n2379) : (n2983 ? (n2379) : (n2976 ? (n2379) : (n2969 ? (n2379) : (n2962 ? (n2379) : (n2955 ? (n2379) : (n2948 ? (n2379) : (n2941 ? (n2379) : (n2934 ? (n2379) : (n2927 ? (n2379) : (n2920 ? (n2379) : (n2913 ? (n2379) : (n2906 ? (n2379) : (n2899 ? (n2379) : (n2892 ? (n2379) : (n2885 ? (n2379) : (n2878 ? (n2379) : (n2871 ? (n2379) : (n2864 ? (n2379) : (n2857 ? (n2379) : (n2850 ? (n2379) : (n2843 ? (n2379) : (n2836 ? (n2379) : (n2829 ? (n2379) : (n2822 ? (n2379) : (n2815 ? (n2379) : (n2808 ? (n2379) : (n2801 ? (n2379) : (n2794 ? (n2379) : (n2787 ? (n2379) : (n2780 ? (n2379) : (n2773 ? (n2379) : (n2766 ? (n2379) : (n2759 ? (n2379) : (n2752 ? (n2379) : (n2745 ? (n2379) : (n2738 ? (n2379) : (n2731 ? (n2379) : (n2724 ? (n2379) : (n2717 ? (n2379) : (n2710 ? (n2379) : (n2703 ? (n2379) : (n2696 ? (n2379) : (n2689 ? (n2379) : (n2682 ? (n2379) : (n2675 ? (n2379) : (n2668 ? (n2379) : (n2661 ? (n2379) : (n2654 ? (n2379) : (n2647 ? (n2379) : (n2640 ? (n2379) : (n2633 ? (n2379) : (n2626 ? (n2379) : (n2619 ? (n2379) : (n2612 ? (n2379) : (n2605 ? (n2379) : (n2598 ? (n2379) : (n2591 ? (n2379) : (n2584 ? (n2379) : (n2577 ? (n2379) : (n2570 ? (n2379) : (n2563 ? (n2379) : (n2556 ? (n2379) : (n2549 ? (n2379) : (n2542 ? (n2379) : (n2535 ? (n2379) : (n2528 ? (n2379) : (n2521 ? (n2379) : (n2514 ? (n2379) : (n2507 ? (n2379) : (n2500 ? (n2379) : (n2493 ? (n2379) : (n2486 ? (n2379) : (n2479 ? (n2379) : (n2472 ? (n2379) : (n2465 ? (n2379) : (n2458 ? (n2379) : (n2451 ? (n2379) : (n2444 ? (n2379) : (n2437 ? (n2379) : (n2430 ? (n2379) : (n2423 ? (n2379) : (n2416 ? (n2379) : (n2409 ? (n2379) : (n2402 ? (n2379) : (n2395 ? (n2379) : (n2388 ? (n2379) : (n2365 ? (n2379) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen6 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_addr7 = n3494 ? (n2380) : (n3487 ? (n2380) : (n3480 ? (n2380) : (n3473 ? (n2380) : (n3466 ? (n2380) : (n3459 ? (n2380) : (n3452 ? (n2380) : (n3445 ? (n2380) : (n3438 ? (n2380) : (n3431 ? (n2380) : (n3424 ? (n2380) : (n3417 ? (n2380) : (n3410 ? (n2380) : (n3403 ? (n2380) : (n3396 ? (n2380) : (n3389 ? (n2380) : (n3382 ? (n2380) : (n3375 ? (n2380) : (n3368 ? (n2380) : (n3361 ? (n2380) : (n3354 ? (n2380) : (n3347 ? (n2380) : (n3340 ? (n2380) : (n3333 ? (n2380) : (n3326 ? (n2380) : (n3319 ? (n2380) : (n3312 ? (n2380) : (n3305 ? (n2380) : (n3298 ? (n2380) : (n3291 ? (n2380) : (n3284 ? (n2380) : (n3277 ? (n2380) : (n3270 ? (n2380) : (n3263 ? (n2380) : (n3256 ? (n2380) : (n3249 ? (n2380) : (n3242 ? (n2380) : (n3235 ? (n2380) : (n3228 ? (n2380) : (n3221 ? (n2380) : (n3214 ? (n2380) : (n3207 ? (n2380) : (n3200 ? (n2380) : (n3193 ? (n2380) : (n3186 ? (n2380) : (n3179 ? (n2380) : (n3172 ? (n2380) : (n3165 ? (n2380) : (n3158 ? (n2380) : (n3151 ? (n2380) : (n3144 ? (n2380) : (n3137 ? (n2380) : (n3130 ? (n2380) : (n3123 ? (n2380) : (n3116 ? (n2380) : (n3109 ? (n2380) : (n3102 ? (n2380) : (n3095 ? (n2380) : (n3088 ? (n2380) : (n3081 ? (n2380) : (n3074 ? (n2380) : (n3067 ? (n2380) : (n3060 ? (n2380) : (n3053 ? (n2380) : (n3046 ? (n2380) : (n3039 ? (n2380) : (n3032 ? (n2380) : (n3025 ? (n2380) : (n3018 ? (n2380) : (n3011 ? (n2380) : (n3004 ? (n2380) : (n2997 ? (n2380) : (n2990 ? (n2380) : (n2983 ? (n2380) : (n2976 ? (n2380) : (n2969 ? (n2380) : (n2962 ? (n2380) : (n2955 ? (n2380) : (n2948 ? (n2380) : (n2941 ? (n2380) : (n2934 ? (n2380) : (n2927 ? (n2380) : (n2920 ? (n2380) : (n2913 ? (n2380) : (n2906 ? (n2380) : (n2899 ? (n2380) : (n2892 ? (n2380) : (n2885 ? (n2380) : (n2878 ? (n2380) : (n2871 ? (n2380) : (n2864 ? (n2380) : (n2857 ? (n2380) : (n2850 ? (n2380) : (n2843 ? (n2380) : (n2836 ? (n2380) : (n2829 ? (n2380) : (n2822 ? (n2380) : (n2815 ? (n2380) : (n2808 ? (n2380) : (n2801 ? (n2380) : (n2794 ? (n2380) : (n2787 ? (n2380) : (n2780 ? (n2380) : (n2773 ? (n2380) : (n2766 ? (n2380) : (n2759 ? (n2380) : (n2752 ? (n2380) : (n2745 ? (n2380) : (n2738 ? (n2380) : (n2731 ? (n2380) : (n2724 ? (n2380) : (n2717 ? (n2380) : (n2710 ? (n2380) : (n2703 ? (n2380) : (n2696 ? (n2380) : (n2689 ? (n2380) : (n2682 ? (n2380) : (n2675 ? (n2380) : (n2668 ? (n2380) : (n2661 ? (n2380) : (n2654 ? (n2380) : (n2647 ? (n2380) : (n2640 ? (n2380) : (n2633 ? (n2380) : (n2626 ? (n2380) : (n2619 ? (n2380) : (n2612 ? (n2380) : (n2605 ? (n2380) : (n2598 ? (n2380) : (n2591 ? (n2380) : (n2584 ? (n2380) : (n2577 ? (n2380) : (n2570 ? (n2380) : (n2563 ? (n2380) : (n2556 ? (n2380) : (n2549 ? (n2380) : (n2542 ? (n2380) : (n2535 ? (n2380) : (n2528 ? (n2380) : (n2521 ? (n2380) : (n2514 ? (n2380) : (n2507 ? (n2380) : (n2500 ? (n2380) : (n2493 ? (n2380) : (n2486 ? (n2380) : (n2479 ? (n2380) : (n2472 ? (n2380) : (n2465 ? (n2380) : (n2458 ? (n2380) : (n2451 ? (n2380) : (n2444 ? (n2380) : (n2437 ? (n2380) : (n2430 ? (n2380) : (n2423 ? (n2380) : (n2416 ? (n2380) : (n2409 ? (n2380) : (n2402 ? (n2380) : (n2395 ? (n2380) : (n2388 ? (n2380) : (n2365 ? (n2380) : (0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_data7 = n3494 ? (n2381) : (n3487 ? (n2381) : (n3480 ? (n2381) : (n3473 ? (n2381) : (n3466 ? (n2381) : (n3459 ? (n2381) : (n3452 ? (n2381) : (n3445 ? (n2381) : (n3438 ? (n2381) : (n3431 ? (n2381) : (n3424 ? (n2381) : (n3417 ? (n2381) : (n3410 ? (n2381) : (n3403 ? (n2381) : (n3396 ? (n2381) : (n3389 ? (n2381) : (n3382 ? (n2381) : (n3375 ? (n2381) : (n3368 ? (n2381) : (n3361 ? (n2381) : (n3354 ? (n2381) : (n3347 ? (n2381) : (n3340 ? (n2381) : (n3333 ? (n2381) : (n3326 ? (n2381) : (n3319 ? (n2381) : (n3312 ? (n2381) : (n3305 ? (n2381) : (n3298 ? (n2381) : (n3291 ? (n2381) : (n3284 ? (n2381) : (n3277 ? (n2381) : (n3270 ? (n2381) : (n3263 ? (n2381) : (n3256 ? (n2381) : (n3249 ? (n2381) : (n3242 ? (n2381) : (n3235 ? (n2381) : (n3228 ? (n2381) : (n3221 ? (n2381) : (n3214 ? (n2381) : (n3207 ? (n2381) : (n3200 ? (n2381) : (n3193 ? (n2381) : (n3186 ? (n2381) : (n3179 ? (n2381) : (n3172 ? (n2381) : (n3165 ? (n2381) : (n3158 ? (n2381) : (n3151 ? (n2381) : (n3144 ? (n2381) : (n3137 ? (n2381) : (n3130 ? (n2381) : (n3123 ? (n2381) : (n3116 ? (n2381) : (n3109 ? (n2381) : (n3102 ? (n2381) : (n3095 ? (n2381) : (n3088 ? (n2381) : (n3081 ? (n2381) : (n3074 ? (n2381) : (n3067 ? (n2381) : (n3060 ? (n2381) : (n3053 ? (n2381) : (n3046 ? (n2381) : (n3039 ? (n2381) : (n3032 ? (n2381) : (n3025 ? (n2381) : (n3018 ? (n2381) : (n3011 ? (n2381) : (n3004 ? (n2381) : (n2997 ? (n2381) : (n2990 ? (n2381) : (n2983 ? (n2381) : (n2976 ? (n2381) : (n2969 ? (n2381) : (n2962 ? (n2381) : (n2955 ? (n2381) : (n2948 ? (n2381) : (n2941 ? (n2381) : (n2934 ? (n2381) : (n2927 ? (n2381) : (n2920 ? (n2381) : (n2913 ? (n2381) : (n2906 ? (n2381) : (n2899 ? (n2381) : (n2892 ? (n2381) : (n2885 ? (n2381) : (n2878 ? (n2381) : (n2871 ? (n2381) : (n2864 ? (n2381) : (n2857 ? (n2381) : (n2850 ? (n2381) : (n2843 ? (n2381) : (n2836 ? (n2381) : (n2829 ? (n2381) : (n2822 ? (n2381) : (n2815 ? (n2381) : (n2808 ? (n2381) : (n2801 ? (n2381) : (n2794 ? (n2381) : (n2787 ? (n2381) : (n2780 ? (n2381) : (n2773 ? (n2381) : (n2766 ? (n2381) : (n2759 ? (n2381) : (n2752 ? (n2381) : (n2745 ? (n2381) : (n2738 ? (n2381) : (n2731 ? (n2381) : (n2724 ? (n2381) : (n2717 ? (n2381) : (n2710 ? (n2381) : (n2703 ? (n2381) : (n2696 ? (n2381) : (n2689 ? (n2381) : (n2682 ? (n2381) : (n2675 ? (n2381) : (n2668 ? (n2381) : (n2661 ? (n2381) : (n2654 ? (n2381) : (n2647 ? (n2381) : (n2640 ? (n2381) : (n2633 ? (n2381) : (n2626 ? (n2381) : (n2619 ? (n2381) : (n2612 ? (n2381) : (n2605 ? (n2381) : (n2598 ? (n2381) : (n2591 ? (n2381) : (n2584 ? (n2381) : (n2577 ? (n2381) : (n2570 ? (n2381) : (n2563 ? (n2381) : (n2556 ? (n2381) : (n2549 ? (n2381) : (n2542 ? (n2381) : (n2535 ? (n2381) : (n2528 ? (n2381) : (n2521 ? (n2381) : (n2514 ? (n2381) : (n2507 ? (n2381) : (n2500 ? (n2381) : (n2493 ? (n2381) : (n2486 ? (n2381) : (n2479 ? (n2381) : (n2472 ? (n2381) : (n2465 ? (n2381) : (n2458 ? (n2381) : (n2451 ? (n2381) : (n2444 ? (n2381) : (n2437 ? (n2381) : (n2430 ? (n2381) : (n2423 ? (n2381) : (n2416 ? (n2381) : (n2409 ? (n2381) : (n2402 ? (n2381) : (n2395 ? (n2381) : (n2388 ? (n2381) : (n2365 ? (n2381) : ('d0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
assign XRAM_wen7 = (n3494) ? ( 1'b1 ) : ((n3487) ? ( 1'b1 ) : ((n3480) ? ( 1'b1 ) : ((n3473) ? ( 1'b1 ) : ((n3466) ? ( 1'b1 ) : ((n3459) ? ( 1'b1 ) : ((n3452) ? ( 1'b1 ) : ((n3445) ? ( 1'b1 ) : ((n3438) ? ( 1'b1 ) : ((n3431) ? ( 1'b1 ) : ((n3424) ? ( 1'b1 ) : ((n3417) ? ( 1'b1 ) : ((n3410) ? ( 1'b1 ) : ((n3403) ? ( 1'b1 ) : ((n3396) ? ( 1'b1 ) : ((n3389) ? ( 1'b1 ) : ((n3382) ? ( 1'b1 ) : ((n3375) ? ( 1'b1 ) : ((n3368) ? ( 1'b1 ) : ((n3361) ? ( 1'b1 ) : ((n3354) ? ( 1'b1 ) : ((n3347) ? ( 1'b1 ) : ((n3340) ? ( 1'b1 ) : ((n3333) ? ( 1'b1 ) : ((n3326) ? ( 1'b1 ) : ((n3319) ? ( 1'b1 ) : ((n3312) ? ( 1'b1 ) : ((n3305) ? ( 1'b1 ) : ((n3298) ? ( 1'b1 ) : ((n3291) ? ( 1'b1 ) : ((n3284) ? ( 1'b1 ) : ((n3277) ? ( 1'b1 ) : ((n3270) ? ( 1'b1 ) : ((n3263) ? ( 1'b1 ) : ((n3256) ? ( 1'b1 ) : ((n3249) ? ( 1'b1 ) : ((n3242) ? ( 1'b1 ) : ((n3235) ? ( 1'b1 ) : ((n3228) ? ( 1'b1 ) : ((n3221) ? ( 1'b1 ) : ((n3214) ? ( 1'b1 ) : ((n3207) ? ( 1'b1 ) : ((n3200) ? ( 1'b1 ) : ((n3193) ? ( 1'b1 ) : ((n3186) ? ( 1'b1 ) : ((n3179) ? ( 1'b1 ) : ((n3172) ? ( 1'b1 ) : ((n3165) ? ( 1'b1 ) : ((n3158) ? ( 1'b1 ) : ((n3151) ? ( 1'b1 ) : ((n3144) ? ( 1'b1 ) : ((n3137) ? ( 1'b1 ) : ((n3130) ? ( 1'b1 ) : ((n3123) ? ( 1'b1 ) : ((n3116) ? ( 1'b1 ) : ((n3109) ? ( 1'b1 ) : ((n3102) ? ( 1'b1 ) : ((n3095) ? ( 1'b1 ) : ((n3088) ? ( 1'b1 ) : ((n3081) ? ( 1'b1 ) : ((n3074) ? ( 1'b1 ) : ((n3067) ? ( 1'b1 ) : ((n3060) ? ( 1'b1 ) : ((n3053) ? ( 1'b1 ) : ((n3046) ? ( 1'b1 ) : ((n3039) ? ( 1'b1 ) : ((n3032) ? ( 1'b1 ) : ((n3025) ? ( 1'b1 ) : ((n3018) ? ( 1'b1 ) : ((n3011) ? ( 1'b1 ) : ((n3004) ? ( 1'b1 ) : ((n2997) ? ( 1'b1 ) : ((n2990) ? ( 1'b1 ) : ((n2983) ? ( 1'b1 ) : ((n2976) ? ( 1'b1 ) : ((n2969) ? ( 1'b1 ) : ((n2962) ? ( 1'b1 ) : ((n2955) ? ( 1'b1 ) : ((n2948) ? ( 1'b1 ) : ((n2941) ? ( 1'b1 ) : ((n2934) ? ( 1'b1 ) : ((n2927) ? ( 1'b1 ) : ((n2920) ? ( 1'b1 ) : ((n2913) ? ( 1'b1 ) : ((n2906) ? ( 1'b1 ) : ((n2899) ? ( 1'b1 ) : ((n2892) ? ( 1'b1 ) : ((n2885) ? ( 1'b1 ) : ((n2878) ? ( 1'b1 ) : ((n2871) ? ( 1'b1 ) : ((n2864) ? ( 1'b1 ) : ((n2857) ? ( 1'b1 ) : ((n2850) ? ( 1'b1 ) : ((n2843) ? ( 1'b1 ) : ((n2836) ? ( 1'b1 ) : ((n2829) ? ( 1'b1 ) : ((n2822) ? ( 1'b1 ) : ((n2815) ? ( 1'b1 ) : ((n2808) ? ( 1'b1 ) : ((n2801) ? ( 1'b1 ) : ((n2794) ? ( 1'b1 ) : ((n2787) ? ( 1'b1 ) : ((n2780) ? ( 1'b1 ) : ((n2773) ? ( 1'b1 ) : ((n2766) ? ( 1'b1 ) : ((n2759) ? ( 1'b1 ) : ((n2752) ? ( 1'b1 ) : ((n2745) ? ( 1'b1 ) : ((n2738) ? ( 1'b1 ) : ((n2731) ? ( 1'b1 ) : ((n2724) ? ( 1'b1 ) : ((n2717) ? ( 1'b1 ) : ((n2710) ? ( 1'b1 ) : ((n2703) ? ( 1'b1 ) : ((n2696) ? ( 1'b1 ) : ((n2689) ? ( 1'b1 ) : ((n2682) ? ( 1'b1 ) : ((n2675) ? ( 1'b1 ) : ((n2668) ? ( 1'b1 ) : ((n2661) ? ( 1'b1 ) : ((n2654) ? ( 1'b1 ) : ((n2647) ? ( 1'b1 ) : ((n2640) ? ( 1'b1 ) : ((n2633) ? ( 1'b1 ) : ((n2626) ? ( 1'b1 ) : ((n2619) ? ( 1'b1 ) : ((n2612) ? ( 1'b1 ) : ((n2605) ? ( 1'b1 ) : ((n2598) ? ( 1'b1 ) : ((n2591) ? ( 1'b1 ) : ((n2584) ? ( 1'b1 ) : ((n2577) ? ( 1'b1 ) : ((n2570) ? ( 1'b1 ) : ((n2563) ? ( 1'b1 ) : ((n2556) ? ( 1'b1 ) : ((n2549) ? ( 1'b1 ) : ((n2542) ? ( 1'b1 ) : ((n2535) ? ( 1'b1 ) : ((n2528) ? ( 1'b1 ) : ((n2521) ? ( 1'b1 ) : ((n2514) ? ( 1'b1 ) : ((n2507) ? ( 1'b1 ) : ((n2500) ? ( 1'b1 ) : ((n2493) ? ( 1'b1 ) : ((n2486) ? ( 1'b1 ) : ((n2479) ? ( 1'b1 ) : ((n2472) ? ( 1'b1 ) : ((n2465) ? ( 1'b1 ) : ((n2458) ? ( 1'b1 ) : ((n2451) ? ( 1'b1 ) : ((n2444) ? ( 1'b1 ) : ((n2437) ? ( 1'b1 ) : ((n2430) ? ( 1'b1 ) : ((n2423) ? ( 1'b1 ) : ((n2416) ? ( 1'b1 ) : ((n2409) ? ( 1'b1 ) : ((n2402) ? ( 1'b1 ) : ((n2395) ? ( 1'b1 ) : ((n2388) ? ( 1'b1 ) : ((n2365) ? ( 1'b1 ) : (1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_sha_valid__) begin
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           dataout <= n649;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           dataout <= n649;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_bytes_read <= n736;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_bytes_read <= n734;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_bytes_read <= n734;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_hs_data <= n824;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_hs_data <= n824;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_len <= n826;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_len <= n828;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_len <= sha_len;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_len <= sha_len;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_rd_data <= n1232;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_rd_data <= n1232;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_rdaddr <= n1234;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_rdaddr <= n1236;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_rdaddr <= sha_rdaddr;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_rdaddr <= sha_rdaddr;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_state <= n1634;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_state <= n1632;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_state <= n1632;
       end
       if ( __ILA_sha_decode_of_I__DOT__0__ && __ILA_sha_grant__[0] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__1__ && __ILA_sha_grant__[1] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__2__ && __ILA_sha_grant__[2] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__3__ && __ILA_sha_grant__[3] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__4__ && __ILA_sha_grant__[4] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__5__ && __ILA_sha_grant__[5] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__6__ && __ILA_sha_grant__[6] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__7__ && __ILA_sha_grant__[7] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__8__ && __ILA_sha_grant__[8] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__9__ && __ILA_sha_grant__[9] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__10__ && __ILA_sha_grant__[10] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__11__ && __ILA_sha_grant__[11] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__12__ && __ILA_sha_grant__[12] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__13__ && __ILA_sha_grant__[13] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__14__ && __ILA_sha_grant__[14] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__15__ && __ILA_sha_grant__[15] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__16__ && __ILA_sha_grant__[16] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__17__ && __ILA_sha_grant__[17] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__18__ && __ILA_sha_grant__[18] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__19__ && __ILA_sha_grant__[19] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__20__ && __ILA_sha_grant__[20] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__21__ && __ILA_sha_grant__[21] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__22__ && __ILA_sha_grant__[22] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__23__ && __ILA_sha_grant__[23] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__24__ && __ILA_sha_grant__[24] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__25__ && __ILA_sha_grant__[25] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__26__ && __ILA_sha_grant__[26] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__27__ && __ILA_sha_grant__[27] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__28__ && __ILA_sha_grant__[28] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__29__ && __ILA_sha_grant__[29] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__30__ && __ILA_sha_grant__[30] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__31__ && __ILA_sha_grant__[31] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__32__ && __ILA_sha_grant__[32] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__33__ && __ILA_sha_grant__[33] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__34__ && __ILA_sha_grant__[34] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__35__ && __ILA_sha_grant__[35] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__36__ && __ILA_sha_grant__[36] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__37__ && __ILA_sha_grant__[37] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__38__ && __ILA_sha_grant__[38] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__39__ && __ILA_sha_grant__[39] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__40__ && __ILA_sha_grant__[40] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__41__ && __ILA_sha_grant__[41] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__42__ && __ILA_sha_grant__[42] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__43__ && __ILA_sha_grant__[43] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__44__ && __ILA_sha_grant__[44] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__45__ && __ILA_sha_grant__[45] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__46__ && __ILA_sha_grant__[46] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__47__ && __ILA_sha_grant__[47] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__48__ && __ILA_sha_grant__[48] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__49__ && __ILA_sha_grant__[49] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__50__ && __ILA_sha_grant__[50] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__51__ && __ILA_sha_grant__[51] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__52__ && __ILA_sha_grant__[52] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__53__ && __ILA_sha_grant__[53] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__54__ && __ILA_sha_grant__[54] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__55__ && __ILA_sha_grant__[55] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__56__ && __ILA_sha_grant__[56] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__57__ && __ILA_sha_grant__[57] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__58__ && __ILA_sha_grant__[58] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__59__ && __ILA_sha_grant__[59] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__60__ && __ILA_sha_grant__[60] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__61__ && __ILA_sha_grant__[61] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__62__ && __ILA_sha_grant__[62] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__63__ && __ILA_sha_grant__[63] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__64__ && __ILA_sha_grant__[64] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__65__ && __ILA_sha_grant__[65] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__66__ && __ILA_sha_grant__[66] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__67__ && __ILA_sha_grant__[67] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__68__ && __ILA_sha_grant__[68] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__69__ && __ILA_sha_grant__[69] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__70__ && __ILA_sha_grant__[70] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__71__ && __ILA_sha_grant__[71] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__72__ && __ILA_sha_grant__[72] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__73__ && __ILA_sha_grant__[73] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__74__ && __ILA_sha_grant__[74] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__75__ && __ILA_sha_grant__[75] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__76__ && __ILA_sha_grant__[76] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__77__ && __ILA_sha_grant__[77] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__78__ && __ILA_sha_grant__[78] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__79__ && __ILA_sha_grant__[79] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__80__ && __ILA_sha_grant__[80] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__81__ && __ILA_sha_grant__[81] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__82__ && __ILA_sha_grant__[82] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__83__ && __ILA_sha_grant__[83] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__84__ && __ILA_sha_grant__[84] ) begin
           sha_wraddr <= n1636;
       end else if ( __ILA_sha_decode_of_I__DOT__85__ && __ILA_sha_grant__[85] ) begin
           sha_wraddr <= n1638;
       end else if ( __ILA_sha_decode_of_I__DOT__86__ && __ILA_sha_grant__[86] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__87__ && __ILA_sha_grant__[87] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__88__ && __ILA_sha_grant__[88] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__89__ && __ILA_sha_grant__[89] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__90__ && __ILA_sha_grant__[90] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__91__ && __ILA_sha_grant__[91] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__92__ && __ILA_sha_grant__[92] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__93__ && __ILA_sha_grant__[93] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__94__ && __ILA_sha_grant__[94] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__95__ && __ILA_sha_grant__[95] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__96__ && __ILA_sha_grant__[96] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__97__ && __ILA_sha_grant__[97] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__98__ && __ILA_sha_grant__[98] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__99__ && __ILA_sha_grant__[99] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__100__ && __ILA_sha_grant__[100] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__101__ && __ILA_sha_grant__[101] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__102__ && __ILA_sha_grant__[102] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__103__ && __ILA_sha_grant__[103] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__104__ && __ILA_sha_grant__[104] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__105__ && __ILA_sha_grant__[105] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__106__ && __ILA_sha_grant__[106] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__107__ && __ILA_sha_grant__[107] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__108__ && __ILA_sha_grant__[108] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__109__ && __ILA_sha_grant__[109] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__110__ && __ILA_sha_grant__[110] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__111__ && __ILA_sha_grant__[111] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__112__ && __ILA_sha_grant__[112] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__113__ && __ILA_sha_grant__[113] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__114__ && __ILA_sha_grant__[114] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__115__ && __ILA_sha_grant__[115] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__116__ && __ILA_sha_grant__[116] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__117__ && __ILA_sha_grant__[117] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__118__ && __ILA_sha_grant__[118] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__119__ && __ILA_sha_grant__[119] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__120__ && __ILA_sha_grant__[120] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__121__ && __ILA_sha_grant__[121] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__122__ && __ILA_sha_grant__[122] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__123__ && __ILA_sha_grant__[123] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__124__ && __ILA_sha_grant__[124] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__125__ && __ILA_sha_grant__[125] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__126__ && __ILA_sha_grant__[126] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__127__ && __ILA_sha_grant__[127] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__128__ && __ILA_sha_grant__[128] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__129__ && __ILA_sha_grant__[129] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__130__ && __ILA_sha_grant__[130] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__131__ && __ILA_sha_grant__[131] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__132__ && __ILA_sha_grant__[132] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__133__ && __ILA_sha_grant__[133] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__134__ && __ILA_sha_grant__[134] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__135__ && __ILA_sha_grant__[135] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__136__ && __ILA_sha_grant__[136] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__137__ && __ILA_sha_grant__[137] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__138__ && __ILA_sha_grant__[138] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__139__ && __ILA_sha_grant__[139] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__140__ && __ILA_sha_grant__[140] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__141__ && __ILA_sha_grant__[141] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__142__ && __ILA_sha_grant__[142] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__143__ && __ILA_sha_grant__[143] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__144__ && __ILA_sha_grant__[144] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__145__ && __ILA_sha_grant__[145] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__146__ && __ILA_sha_grant__[146] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__147__ && __ILA_sha_grant__[147] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__148__ && __ILA_sha_grant__[148] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__149__ && __ILA_sha_grant__[149] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__150__ && __ILA_sha_grant__[150] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__151__ && __ILA_sha_grant__[151] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__152__ && __ILA_sha_grant__[152] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__153__ && __ILA_sha_grant__[153] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__154__ && __ILA_sha_grant__[154] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__155__ && __ILA_sha_grant__[155] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__156__ && __ILA_sha_grant__[156] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__157__ && __ILA_sha_grant__[157] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__158__ && __ILA_sha_grant__[158] ) begin
           sha_wraddr <= sha_wraddr;
       end else if ( __ILA_sha_decode_of_I__DOT__159__ && __ILA_sha_grant__[159] ) begin
           sha_wraddr <= sha_wraddr;
       end
   end
end
endmodule
