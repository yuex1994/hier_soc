module AES(
__ILA_AES_grant__,
clk,
cmd,
cmdaddr,
cmddata,
nondet_unknown0_n72,
nondet_unknown1_n75,
nondet_unknown2_n175,
rst,
__ILA_AES_acc_decode__,
__ILA_AES_decode_of_GET_STATUS__,
__ILA_AES_decode_of_READ_ADDRESS__,
__ILA_AES_decode_of_READ_COUNTER__,
__ILA_AES_decode_of_READ_KEY__,
__ILA_AES_decode_of_READ_LENGTH__,
__ILA_AES_decode_of_START_ENCRYPT__,
__ILA_AES_decode_of_WRITE_ADDRESS__,
__ILA_AES_decode_of_WRITE_COUNTER__,
__ILA_AES_decode_of_WRITE_KEY__,
__ILA_AES_decode_of_WRITE_LENGTH__,
__ILA_AES_valid__,
aes_status,
aes_address,
aes_length,
aes_counter,
aes_key,
outdata
);
input      [9:0] __ILA_AES_grant__;
input            clk;
input      [1:0] cmd;
input     [15:0] cmdaddr;
input      [7:0] cmddata;
input      [1:0] nondet_unknown0_n72;
input      [1:0] nondet_unknown1_n75;
input    [127:0] nondet_unknown2_n175;
input            rst;
output      [9:0] __ILA_AES_acc_decode__;
output            __ILA_AES_decode_of_GET_STATUS__;
output            __ILA_AES_decode_of_READ_ADDRESS__;
output            __ILA_AES_decode_of_READ_COUNTER__;
output            __ILA_AES_decode_of_READ_KEY__;
output            __ILA_AES_decode_of_READ_LENGTH__;
output            __ILA_AES_decode_of_START_ENCRYPT__;
output            __ILA_AES_decode_of_WRITE_ADDRESS__;
output            __ILA_AES_decode_of_WRITE_COUNTER__;
output            __ILA_AES_decode_of_WRITE_KEY__;
output            __ILA_AES_decode_of_WRITE_LENGTH__;
output            __ILA_AES_valid__;
output reg      [1:0] aes_status;
output reg     [15:0] aes_address;
output reg     [15:0] aes_length;
output reg    [127:0] aes_counter;
output reg    [127:0] aes_key;
output reg      [7:0] outdata;
wire      [9:0] __ILA_AES_acc_decode__;
wire            __ILA_AES_decode_of_GET_STATUS__;
wire            __ILA_AES_decode_of_READ_ADDRESS__;
wire            __ILA_AES_decode_of_READ_COUNTER__;
wire            __ILA_AES_decode_of_READ_KEY__;
wire            __ILA_AES_decode_of_READ_LENGTH__;
wire            __ILA_AES_decode_of_START_ENCRYPT__;
wire            __ILA_AES_decode_of_WRITE_ADDRESS__;
wire            __ILA_AES_decode_of_WRITE_COUNTER__;
wire            __ILA_AES_decode_of_WRITE_KEY__;
wire            __ILA_AES_decode_of_WRITE_LENGTH__;
wire      [9:0] __ILA_AES_grant__;
wire            __ILA_AES_valid__;
wire            clk;
wire      [1:0] cmd;
wire     [15:0] cmdaddr;
wire      [7:0] cmddata;
wire            n0;
wire            n1;
wire            n10;
wire     [15:0] n100;
wire            n101;
wire      [7:0] n102;
wire      [7:0] n103;
wire     [15:0] n104;
wire            n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire     [15:0] n108;
wire            n109;
wire            n11;
wire      [7:0] n110;
wire      [7:0] n111;
wire     [15:0] n112;
wire            n113;
wire      [7:0] n114;
wire      [7:0] n115;
wire     [15:0] n116;
wire            n117;
wire      [7:0] n118;
wire      [7:0] n119;
wire            n12;
wire     [15:0] n120;
wire            n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire     [15:0] n124;
wire            n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire     [15:0] n128;
wire            n129;
wire            n13;
wire      [7:0] n130;
wire      [7:0] n131;
wire     [15:0] n132;
wire            n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire     [15:0] n136;
wire            n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire            n14;
wire     [15:0] n140;
wire            n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire     [15:0] n144;
wire            n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire     [15:0] n148;
wire            n149;
wire            n15;
wire      [7:0] n150;
wire      [7:0] n151;
wire     [15:0] n152;
wire            n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire     [15:0] n156;
wire            n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire            n16;
wire     [15:0] n160;
wire     [23:0] n161;
wire     [31:0] n162;
wire     [39:0] n163;
wire     [47:0] n164;
wire     [55:0] n165;
wire     [63:0] n166;
wire     [71:0] n167;
wire     [79:0] n168;
wire     [87:0] n169;
wire            n17;
wire     [95:0] n170;
wire    [103:0] n171;
wire    [111:0] n172;
wire    [119:0] n173;
wire    [127:0] n174;
wire    [127:0] n176;
wire    [127:0] n177;
wire     [15:0] n178;
wire            n179;
wire            n18;
wire      [7:0] n180;
wire      [7:0] n181;
wire     [15:0] n182;
wire            n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire     [15:0] n186;
wire            n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire            n19;
wire     [15:0] n190;
wire            n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire     [15:0] n194;
wire            n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire     [15:0] n198;
wire            n199;
wire            n2;
wire            n20;
wire      [7:0] n200;
wire      [7:0] n201;
wire     [15:0] n202;
wire            n203;
wire      [7:0] n204;
wire      [7:0] n205;
wire     [15:0] n206;
wire            n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire            n21;
wire     [15:0] n210;
wire            n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire     [15:0] n214;
wire            n215;
wire      [7:0] n216;
wire      [7:0] n217;
wire     [15:0] n218;
wire            n219;
wire            n22;
wire      [7:0] n220;
wire      [7:0] n221;
wire     [15:0] n222;
wire            n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire     [15:0] n226;
wire            n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire            n23;
wire     [15:0] n230;
wire            n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire     [15:0] n234;
wire            n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire     [15:0] n238;
wire            n239;
wire            n24;
wire      [7:0] n240;
wire      [7:0] n241;
wire     [15:0] n242;
wire     [23:0] n243;
wire     [31:0] n244;
wire     [39:0] n245;
wire     [47:0] n246;
wire     [55:0] n247;
wire     [63:0] n248;
wire     [71:0] n249;
wire            n25;
wire     [79:0] n250;
wire     [87:0] n251;
wire     [95:0] n252;
wire    [103:0] n253;
wire    [111:0] n254;
wire    [119:0] n255;
wire    [127:0] n256;
wire    [127:0] n257;
wire     [15:0] n258;
wire            n259;
wire            n26;
wire      [7:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire     [15:0] n263;
wire            n264;
wire      [7:0] n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire     [15:0] n268;
wire            n269;
wire            n27;
wire      [7:0] n270;
wire     [15:0] n271;
wire            n272;
wire      [7:0] n273;
wire     [15:0] n274;
wire            n275;
wire      [7:0] n276;
wire     [15:0] n277;
wire            n278;
wire      [7:0] n279;
wire            n28;
wire     [15:0] n280;
wire            n281;
wire      [7:0] n282;
wire     [15:0] n283;
wire            n284;
wire      [7:0] n285;
wire     [15:0] n286;
wire            n287;
wire      [7:0] n288;
wire     [15:0] n289;
wire            n29;
wire            n290;
wire      [7:0] n291;
wire     [15:0] n292;
wire            n293;
wire      [7:0] n294;
wire     [15:0] n295;
wire            n296;
wire      [7:0] n297;
wire     [15:0] n298;
wire            n299;
wire            n3;
wire            n30;
wire      [7:0] n300;
wire     [15:0] n301;
wire            n302;
wire      [7:0] n303;
wire     [15:0] n304;
wire            n305;
wire      [7:0] n306;
wire     [15:0] n307;
wire            n308;
wire      [7:0] n309;
wire            n31;
wire     [15:0] n310;
wire            n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire            n32;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire     [15:0] n329;
wire            n33;
wire            n330;
wire      [7:0] n331;
wire     [15:0] n332;
wire            n333;
wire      [7:0] n334;
wire     [15:0] n335;
wire            n336;
wire      [7:0] n337;
wire     [15:0] n338;
wire            n339;
wire            n34;
wire      [7:0] n340;
wire     [15:0] n341;
wire            n342;
wire      [7:0] n343;
wire     [15:0] n344;
wire            n345;
wire      [7:0] n346;
wire     [15:0] n347;
wire            n348;
wire      [7:0] n349;
wire            n35;
wire     [15:0] n350;
wire            n351;
wire      [7:0] n352;
wire     [15:0] n353;
wire            n354;
wire      [7:0] n355;
wire     [15:0] n356;
wire            n357;
wire      [7:0] n358;
wire     [15:0] n359;
wire            n36;
wire            n360;
wire      [7:0] n361;
wire     [15:0] n362;
wire            n363;
wire      [7:0] n364;
wire     [15:0] n365;
wire            n366;
wire      [7:0] n367;
wire     [15:0] n368;
wire            n369;
wire            n37;
wire      [7:0] n370;
wire     [15:0] n371;
wire            n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire            n38;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire            n39;
wire     [15:0] n390;
wire            n391;
wire      [7:0] n392;
wire     [15:0] n393;
wire            n394;
wire      [7:0] n395;
wire     [15:0] n396;
wire            n397;
wire      [7:0] n398;
wire     [15:0] n399;
wire            n4;
wire            n40;
wire            n400;
wire      [7:0] n401;
wire     [15:0] n402;
wire            n403;
wire      [7:0] n404;
wire     [15:0] n405;
wire            n406;
wire      [7:0] n407;
wire     [15:0] n408;
wire            n409;
wire            n41;
wire      [7:0] n410;
wire     [15:0] n411;
wire            n412;
wire      [7:0] n413;
wire     [15:0] n414;
wire            n415;
wire      [7:0] n416;
wire     [15:0] n417;
wire            n418;
wire      [7:0] n419;
wire            n42;
wire     [15:0] n420;
wire            n421;
wire      [7:0] n422;
wire     [15:0] n423;
wire            n424;
wire      [7:0] n425;
wire     [15:0] n426;
wire            n427;
wire      [7:0] n428;
wire     [15:0] n429;
wire            n43;
wire            n430;
wire      [7:0] n431;
wire     [15:0] n432;
wire            n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire            n44;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire            n45;
wire      [7:0] n450;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire            n5;
wire            n50;
wire            n51;
wire            n52;
wire            n53;
wire            n54;
wire            n55;
wire            n56;
wire            n57;
wire            n58;
wire            n59;
wire            n6;
wire            n60;
wire            n61;
wire            n62;
wire            n63;
wire            n64;
wire            n65;
wire            n66;
wire            n67;
wire            n68;
wire            n69;
wire            n7;
wire            n70;
wire            n71;
wire      [1:0] n73;
wire      [1:0] n74;
wire      [1:0] n76;
wire      [1:0] n77;
wire            n78;
wire      [7:0] n79;
wire            n8;
wire      [7:0] n80;
wire            n81;
wire      [7:0] n82;
wire      [7:0] n83;
wire     [15:0] n84;
wire     [15:0] n85;
wire     [15:0] n86;
wire            n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire            n9;
wire     [15:0] n90;
wire            n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire     [15:0] n94;
wire     [15:0] n95;
wire     [15:0] n96;
wire            n97;
wire      [7:0] n98;
wire      [7:0] n99;
wire      [1:0] nondet_unknown0_n72;
wire      [1:0] nondet_unknown1_n75;
wire    [127:0] nondet_unknown2_n175;
wire            rst;
assign n0 =  ( cmd ) == ( 2'd1 )  ;
assign n1 =  ( cmd ) == ( 2'd2 )  ;
assign n2 =  ( n0 ) | ( n1 )  ;
assign __ILA_AES_valid__ = n2 ;
assign n3 =  ( cmd ) == ( 2'd2 )  ;
assign n4 =  ( cmdaddr ) == ( 16'd65282 )  ;
assign n5 =  ( cmdaddr ) > ( 16'd65282 )  ;
assign n6 =  ( n4 ) | ( n5 )  ;
assign n7 =  ( n3 ) & (n6 )  ;
assign n8 =  ( cmdaddr ) < ( 16'd65284 )  ;
assign n9 =  ( n7 ) & (n8 )  ;
assign __ILA_AES_decode_of_WRITE_ADDRESS__ = n9 ;
assign __ILA_AES_acc_decode__[0] = __ILA_AES_decode_of_WRITE_ADDRESS__ ;
assign n10 =  ( cmd ) == ( 2'd2 )  ;
assign n11 =  ( cmdaddr ) == ( 16'd65280 )  ;
assign n12 =  ( n10 ) & (n11 )  ;
assign n13 =  ( cmddata ) == ( 8'd1 )  ;
assign n14 =  ( n12 ) & (n13 )  ;
assign __ILA_AES_decode_of_START_ENCRYPT__ = n14 ;
assign __ILA_AES_acc_decode__[1] = __ILA_AES_decode_of_START_ENCRYPT__ ;
assign n15 =  ( cmd ) == ( 2'd1 )  ;
assign n16 =  ( cmdaddr ) == ( 16'd65284 )  ;
assign n17 =  ( cmdaddr ) > ( 16'd65284 )  ;
assign n18 =  ( n16 ) | ( n17 )  ;
assign n19 =  ( n15 ) & (n18 )  ;
assign n20 =  ( cmdaddr ) < ( 16'd65286 )  ;
assign n21 =  ( n19 ) & (n20 )  ;
assign __ILA_AES_decode_of_READ_LENGTH__ = n21 ;
assign __ILA_AES_acc_decode__[2] = __ILA_AES_decode_of_READ_LENGTH__ ;
assign n22 =  ( cmd ) == ( 2'd1 )  ;
assign n23 =  ( cmdaddr ) == ( 16'd65282 )  ;
assign n24 =  ( cmdaddr ) > ( 16'd65282 )  ;
assign n25 =  ( n23 ) | ( n24 )  ;
assign n26 =  ( n22 ) & (n25 )  ;
assign n27 =  ( cmdaddr ) < ( 16'd65284 )  ;
assign n28 =  ( n26 ) & (n27 )  ;
assign __ILA_AES_decode_of_READ_ADDRESS__ = n28 ;
assign __ILA_AES_acc_decode__[3] = __ILA_AES_decode_of_READ_ADDRESS__ ;
assign n29 =  ( cmd ) == ( 2'd1 )  ;
assign n30 =  ( cmdaddr ) == ( 16'd65312 )  ;
assign n31 =  ( cmdaddr ) > ( 16'd65312 )  ;
assign n32 =  ( n30 ) | ( n31 )  ;
assign n33 =  ( n29 ) & (n32 )  ;
assign n34 =  ( cmdaddr ) < ( 16'd65328 )  ;
assign n35 =  ( n33 ) & (n34 )  ;
assign __ILA_AES_decode_of_READ_KEY__ = n35 ;
assign __ILA_AES_acc_decode__[4] = __ILA_AES_decode_of_READ_KEY__ ;
assign n36 =  ( cmd ) == ( 2'd1 )  ;
assign n37 =  ( cmdaddr ) == ( 16'd65296 )  ;
assign n38 =  ( cmdaddr ) > ( 16'd65296 )  ;
assign n39 =  ( n37 ) | ( n38 )  ;
assign n40 =  ( n36 ) & (n39 )  ;
assign n41 =  ( cmdaddr ) < ( 16'd65312 )  ;
assign n42 =  ( n40 ) & (n41 )  ;
assign __ILA_AES_decode_of_READ_COUNTER__ = n42 ;
assign __ILA_AES_acc_decode__[5] = __ILA_AES_decode_of_READ_COUNTER__ ;
assign n43 =  ( cmd ) == ( 2'd1 )  ;
assign n44 =  ( cmdaddr ) == ( 16'd65296 )  ;
assign n45 =  ( cmdaddr ) > ( 16'd65296 )  ;
assign n46 =  ( n44 ) | ( n45 )  ;
assign n47 =  ( n43 ) & (n46 )  ;
assign n48 =  ( cmdaddr ) < ( 16'd65312 )  ;
assign n49 =  ( n47 ) & (n48 )  ;
assign __ILA_AES_decode_of_GET_STATUS__ = n49 ;
assign __ILA_AES_acc_decode__[6] = __ILA_AES_decode_of_GET_STATUS__ ;
assign n50 =  ( cmd ) == ( 2'd2 )  ;
assign n51 =  ( cmdaddr ) == ( 16'd65284 )  ;
assign n52 =  ( cmdaddr ) > ( 16'd65284 )  ;
assign n53 =  ( n51 ) | ( n52 )  ;
assign n54 =  ( n50 ) & (n53 )  ;
assign n55 =  ( cmdaddr ) < ( 16'd65286 )  ;
assign n56 =  ( n54 ) & (n55 )  ;
assign __ILA_AES_decode_of_WRITE_LENGTH__ = n56 ;
assign __ILA_AES_acc_decode__[7] = __ILA_AES_decode_of_WRITE_LENGTH__ ;
assign n57 =  ( cmd ) == ( 2'd2 )  ;
assign n58 =  ( cmdaddr ) == ( 16'd65312 )  ;
assign n59 =  ( cmdaddr ) > ( 16'd65312 )  ;
assign n60 =  ( n58 ) | ( n59 )  ;
assign n61 =  ( n57 ) & (n60 )  ;
assign n62 =  ( cmdaddr ) < ( 16'd65328 )  ;
assign n63 =  ( n61 ) & (n62 )  ;
assign __ILA_AES_decode_of_WRITE_KEY__ = n63 ;
assign __ILA_AES_acc_decode__[8] = __ILA_AES_decode_of_WRITE_KEY__ ;
assign n64 =  ( cmd ) == ( 2'd2 )  ;
assign n65 =  ( cmdaddr ) == ( 16'd65296 )  ;
assign n66 =  ( cmdaddr ) > ( 16'd65296 )  ;
assign n67 =  ( n65 ) | ( n66 )  ;
assign n68 =  ( n64 ) & (n67 )  ;
assign n69 =  ( cmdaddr ) < ( 16'd65312 )  ;
assign n70 =  ( n68 ) & (n69 )  ;
assign __ILA_AES_decode_of_WRITE_COUNTER__ = n70 ;
assign __ILA_AES_acc_decode__[9] = __ILA_AES_decode_of_WRITE_COUNTER__ ;
assign n71 =  ( aes_status ) == ( 2'd0 )  ;
assign n73 = nondet_unknown0_n72 ;
assign n74 =  ( n71 ) ? ( 2'd1 ) : ( n73 ) ;
assign n76 = nondet_unknown1_n75 ;
assign n77 =  ( n71 ) ? ( aes_status ) : ( n76 ) ;
assign n78 =  ( cmdaddr ) == ( 16'd65283 )  ;
assign n79 = aes_address[15:8] ;
assign n80 =  ( n78 ) ? ( cmddata ) : ( n79 ) ;
assign n81 =  ( cmdaddr ) == ( 16'd65282 )  ;
assign n82 = aes_address[7:0] ;
assign n83 =  ( n81 ) ? ( cmddata ) : ( n82 ) ;
assign n84 =  { ( n80 ) , ( n83 ) }  ;
assign n85 =  ( n71 ) ? ( n84 ) : ( aes_address ) ;
assign n86 =  ( cmdaddr ) - ( 16'd65284 )  ;
assign n87 =  ( n86 ) == ( 16'd1 )  ;
assign n88 = aes_length[15:8] ;
assign n89 =  ( n87 ) ? ( cmddata ) : ( n88 ) ;
assign n90 =  ( cmdaddr ) - ( 16'd65284 )  ;
assign n91 =  ( n90 ) == ( 16'd0 )  ;
assign n92 = aes_length[7:0] ;
assign n93 =  ( n91 ) ? ( cmddata ) : ( n92 ) ;
assign n94 =  { ( n89 ) , ( n93 ) }  ;
assign n95 =  ( n71 ) ? ( n94 ) : ( aes_length ) ;
assign n96 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n97 =  ( n96 ) == ( 16'd15 )  ;
assign n98 = aes_counter[127:120] ;
assign n99 =  ( n97 ) ? ( cmddata ) : ( n98 ) ;
assign n100 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n101 =  ( n100 ) == ( 16'd14 )  ;
assign n102 = aes_counter[119:112] ;
assign n103 =  ( n101 ) ? ( cmddata ) : ( n102 ) ;
assign n104 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n105 =  ( n104 ) == ( 16'd13 )  ;
assign n106 = aes_counter[111:104] ;
assign n107 =  ( n105 ) ? ( cmddata ) : ( n106 ) ;
assign n108 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n109 =  ( n108 ) == ( 16'd12 )  ;
assign n110 = aes_counter[103:96] ;
assign n111 =  ( n109 ) ? ( cmddata ) : ( n110 ) ;
assign n112 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n113 =  ( n112 ) == ( 16'd11 )  ;
assign n114 = aes_counter[95:88] ;
assign n115 =  ( n113 ) ? ( cmddata ) : ( n114 ) ;
assign n116 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n117 =  ( n116 ) == ( 16'd10 )  ;
assign n118 = aes_counter[87:80] ;
assign n119 =  ( n117 ) ? ( cmddata ) : ( n118 ) ;
assign n120 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n121 =  ( n120 ) == ( 16'd9 )  ;
assign n122 = aes_counter[79:72] ;
assign n123 =  ( n121 ) ? ( cmddata ) : ( n122 ) ;
assign n124 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n125 =  ( n124 ) == ( 16'd8 )  ;
assign n126 = aes_counter[71:64] ;
assign n127 =  ( n125 ) ? ( cmddata ) : ( n126 ) ;
assign n128 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n129 =  ( n128 ) == ( 16'd7 )  ;
assign n130 = aes_counter[63:56] ;
assign n131 =  ( n129 ) ? ( cmddata ) : ( n130 ) ;
assign n132 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n133 =  ( n132 ) == ( 16'd6 )  ;
assign n134 = aes_counter[55:48] ;
assign n135 =  ( n133 ) ? ( cmddata ) : ( n134 ) ;
assign n136 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n137 =  ( n136 ) == ( 16'd5 )  ;
assign n138 = aes_counter[47:40] ;
assign n139 =  ( n137 ) ? ( cmddata ) : ( n138 ) ;
assign n140 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n141 =  ( n140 ) == ( 16'd4 )  ;
assign n142 = aes_counter[39:32] ;
assign n143 =  ( n141 ) ? ( cmddata ) : ( n142 ) ;
assign n144 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n145 =  ( n144 ) == ( 16'd3 )  ;
assign n146 = aes_counter[31:24] ;
assign n147 =  ( n145 ) ? ( cmddata ) : ( n146 ) ;
assign n148 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n149 =  ( n148 ) == ( 16'd2 )  ;
assign n150 = aes_counter[23:16] ;
assign n151 =  ( n149 ) ? ( cmddata ) : ( n150 ) ;
assign n152 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n153 =  ( n152 ) == ( 16'd1 )  ;
assign n154 = aes_counter[15:8] ;
assign n155 =  ( n153 ) ? ( cmddata ) : ( n154 ) ;
assign n156 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n157 =  ( n156 ) == ( 16'd0 )  ;
assign n158 = aes_counter[7:0] ;
assign n159 =  ( n157 ) ? ( cmddata ) : ( n158 ) ;
assign n160 =  { ( n155 ) , ( n159 ) }  ;
assign n161 =  { ( n151 ) , ( n160 ) }  ;
assign n162 =  { ( n147 ) , ( n161 ) }  ;
assign n163 =  { ( n143 ) , ( n162 ) }  ;
assign n164 =  { ( n139 ) , ( n163 ) }  ;
assign n165 =  { ( n135 ) , ( n164 ) }  ;
assign n166 =  { ( n131 ) , ( n165 ) }  ;
assign n167 =  { ( n127 ) , ( n166 ) }  ;
assign n168 =  { ( n123 ) , ( n167 ) }  ;
assign n169 =  { ( n119 ) , ( n168 ) }  ;
assign n170 =  { ( n115 ) , ( n169 ) }  ;
assign n171 =  { ( n111 ) , ( n170 ) }  ;
assign n172 =  { ( n107 ) , ( n171 ) }  ;
assign n173 =  { ( n103 ) , ( n172 ) }  ;
assign n174 =  { ( n99 ) , ( n173 ) }  ;
assign n176 = nondet_unknown2_n175 ;
assign n177 =  ( n71 ) ? ( n174 ) : ( n176 ) ;
assign n178 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n179 =  ( n178 ) == ( 16'd15 )  ;
assign n180 = aes_key[127:120] ;
assign n181 =  ( n179 ) ? ( cmddata ) : ( n180 ) ;
assign n182 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n183 =  ( n182 ) == ( 16'd14 )  ;
assign n184 = aes_key[119:112] ;
assign n185 =  ( n183 ) ? ( cmddata ) : ( n184 ) ;
assign n186 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n187 =  ( n186 ) == ( 16'd13 )  ;
assign n188 = aes_key[111:104] ;
assign n189 =  ( n187 ) ? ( cmddata ) : ( n188 ) ;
assign n190 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n191 =  ( n190 ) == ( 16'd12 )  ;
assign n192 = aes_key[103:96] ;
assign n193 =  ( n191 ) ? ( cmddata ) : ( n192 ) ;
assign n194 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n195 =  ( n194 ) == ( 16'd11 )  ;
assign n196 = aes_key[95:88] ;
assign n197 =  ( n195 ) ? ( cmddata ) : ( n196 ) ;
assign n198 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n199 =  ( n198 ) == ( 16'd10 )  ;
assign n200 = aes_key[87:80] ;
assign n201 =  ( n199 ) ? ( cmddata ) : ( n200 ) ;
assign n202 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n203 =  ( n202 ) == ( 16'd9 )  ;
assign n204 = aes_key[79:72] ;
assign n205 =  ( n203 ) ? ( cmddata ) : ( n204 ) ;
assign n206 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n207 =  ( n206 ) == ( 16'd8 )  ;
assign n208 = aes_key[71:64] ;
assign n209 =  ( n207 ) ? ( cmddata ) : ( n208 ) ;
assign n210 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n211 =  ( n210 ) == ( 16'd7 )  ;
assign n212 = aes_key[63:56] ;
assign n213 =  ( n211 ) ? ( cmddata ) : ( n212 ) ;
assign n214 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n215 =  ( n214 ) == ( 16'd6 )  ;
assign n216 = aes_key[55:48] ;
assign n217 =  ( n215 ) ? ( cmddata ) : ( n216 ) ;
assign n218 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n219 =  ( n218 ) == ( 16'd5 )  ;
assign n220 = aes_key[47:40] ;
assign n221 =  ( n219 ) ? ( cmddata ) : ( n220 ) ;
assign n222 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n223 =  ( n222 ) == ( 16'd4 )  ;
assign n224 = aes_key[39:32] ;
assign n225 =  ( n223 ) ? ( cmddata ) : ( n224 ) ;
assign n226 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n227 =  ( n226 ) == ( 16'd3 )  ;
assign n228 = aes_key[31:24] ;
assign n229 =  ( n227 ) ? ( cmddata ) : ( n228 ) ;
assign n230 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n231 =  ( n230 ) == ( 16'd2 )  ;
assign n232 = aes_key[23:16] ;
assign n233 =  ( n231 ) ? ( cmddata ) : ( n232 ) ;
assign n234 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n235 =  ( n234 ) == ( 16'd1 )  ;
assign n236 = aes_key[15:8] ;
assign n237 =  ( n235 ) ? ( cmddata ) : ( n236 ) ;
assign n238 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n239 =  ( n238 ) == ( 16'd0 )  ;
assign n240 = aes_key[7:0] ;
assign n241 =  ( n239 ) ? ( cmddata ) : ( n240 ) ;
assign n242 =  { ( n237 ) , ( n241 ) }  ;
assign n243 =  { ( n233 ) , ( n242 ) }  ;
assign n244 =  { ( n229 ) , ( n243 ) }  ;
assign n245 =  { ( n225 ) , ( n244 ) }  ;
assign n246 =  { ( n221 ) , ( n245 ) }  ;
assign n247 =  { ( n217 ) , ( n246 ) }  ;
assign n248 =  { ( n213 ) , ( n247 ) }  ;
assign n249 =  { ( n209 ) , ( n248 ) }  ;
assign n250 =  { ( n205 ) , ( n249 ) }  ;
assign n251 =  { ( n201 ) , ( n250 ) }  ;
assign n252 =  { ( n197 ) , ( n251 ) }  ;
assign n253 =  { ( n193 ) , ( n252 ) }  ;
assign n254 =  { ( n189 ) , ( n253 ) }  ;
assign n255 =  { ( n185 ) , ( n254 ) }  ;
assign n256 =  { ( n181 ) , ( n255 ) }  ;
assign n257 =  ( n71 ) ? ( n256 ) : ( aes_key ) ;
assign n258 =  ( cmdaddr ) - ( 16'd65284 )  ;
assign n259 =  ( n258 ) == ( 16'd1 )  ;
assign n260 = aes_length[15:8] ;
assign n261 = aes_length[7:0] ;
assign n262 =  ( n259 ) ? ( n260 ) : ( n261 ) ;
assign n263 =  ( cmdaddr ) - ( 16'd65282 )  ;
assign n264 =  ( n263 ) == ( 16'd1 )  ;
assign n265 = aes_address[15:8] ;
assign n266 = aes_address[7:0] ;
assign n267 =  ( n264 ) ? ( n265 ) : ( n266 ) ;
assign n268 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n269 =  ( n268 ) == ( 16'd15 )  ;
assign n270 = aes_key[127:120] ;
assign n271 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n272 =  ( n271 ) == ( 16'd14 )  ;
assign n273 = aes_key[119:112] ;
assign n274 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n275 =  ( n274 ) == ( 16'd13 )  ;
assign n276 = aes_key[111:104] ;
assign n277 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n278 =  ( n277 ) == ( 16'd12 )  ;
assign n279 = aes_key[103:96] ;
assign n280 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n281 =  ( n280 ) == ( 16'd11 )  ;
assign n282 = aes_key[95:88] ;
assign n283 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n284 =  ( n283 ) == ( 16'd10 )  ;
assign n285 = aes_key[87:80] ;
assign n286 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n287 =  ( n286 ) == ( 16'd9 )  ;
assign n288 = aes_key[79:72] ;
assign n289 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n290 =  ( n289 ) == ( 16'd8 )  ;
assign n291 = aes_key[71:64] ;
assign n292 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n293 =  ( n292 ) == ( 16'd7 )  ;
assign n294 = aes_key[63:56] ;
assign n295 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n296 =  ( n295 ) == ( 16'd6 )  ;
assign n297 = aes_key[55:48] ;
assign n298 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n299 =  ( n298 ) == ( 16'd5 )  ;
assign n300 = aes_key[47:40] ;
assign n301 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n302 =  ( n301 ) == ( 16'd4 )  ;
assign n303 = aes_key[39:32] ;
assign n304 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n305 =  ( n304 ) == ( 16'd3 )  ;
assign n306 = aes_key[31:24] ;
assign n307 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n308 =  ( n307 ) == ( 16'd2 )  ;
assign n309 = aes_key[23:16] ;
assign n310 =  ( cmdaddr ) - ( 16'd65312 )  ;
assign n311 =  ( n310 ) == ( 16'd1 )  ;
assign n312 = aes_key[15:8] ;
assign n313 = aes_key[7:0] ;
assign n314 =  ( n311 ) ? ( n312 ) : ( n313 ) ;
assign n315 =  ( n308 ) ? ( n309 ) : ( n314 ) ;
assign n316 =  ( n305 ) ? ( n306 ) : ( n315 ) ;
assign n317 =  ( n302 ) ? ( n303 ) : ( n316 ) ;
assign n318 =  ( n299 ) ? ( n300 ) : ( n317 ) ;
assign n319 =  ( n296 ) ? ( n297 ) : ( n318 ) ;
assign n320 =  ( n293 ) ? ( n294 ) : ( n319 ) ;
assign n321 =  ( n290 ) ? ( n291 ) : ( n320 ) ;
assign n322 =  ( n287 ) ? ( n288 ) : ( n321 ) ;
assign n323 =  ( n284 ) ? ( n285 ) : ( n322 ) ;
assign n324 =  ( n281 ) ? ( n282 ) : ( n323 ) ;
assign n325 =  ( n278 ) ? ( n279 ) : ( n324 ) ;
assign n326 =  ( n275 ) ? ( n276 ) : ( n325 ) ;
assign n327 =  ( n272 ) ? ( n273 ) : ( n326 ) ;
assign n328 =  ( n269 ) ? ( n270 ) : ( n327 ) ;
assign n329 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n330 =  ( n329 ) == ( 16'd15 )  ;
assign n331 = aes_counter[127:120] ;
assign n332 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n333 =  ( n332 ) == ( 16'd14 )  ;
assign n334 = aes_counter[119:112] ;
assign n335 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n336 =  ( n335 ) == ( 16'd13 )  ;
assign n337 = aes_counter[111:104] ;
assign n338 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n339 =  ( n338 ) == ( 16'd12 )  ;
assign n340 = aes_counter[103:96] ;
assign n341 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n342 =  ( n341 ) == ( 16'd11 )  ;
assign n343 = aes_counter[95:88] ;
assign n344 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n345 =  ( n344 ) == ( 16'd10 )  ;
assign n346 = aes_counter[87:80] ;
assign n347 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n348 =  ( n347 ) == ( 16'd9 )  ;
assign n349 = aes_counter[79:72] ;
assign n350 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n351 =  ( n350 ) == ( 16'd8 )  ;
assign n352 = aes_counter[71:64] ;
assign n353 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n354 =  ( n353 ) == ( 16'd7 )  ;
assign n355 = aes_counter[63:56] ;
assign n356 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n357 =  ( n356 ) == ( 16'd6 )  ;
assign n358 = aes_counter[55:48] ;
assign n359 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n360 =  ( n359 ) == ( 16'd5 )  ;
assign n361 = aes_counter[47:40] ;
assign n362 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n363 =  ( n362 ) == ( 16'd4 )  ;
assign n364 = aes_counter[39:32] ;
assign n365 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n366 =  ( n365 ) == ( 16'd3 )  ;
assign n367 = aes_counter[31:24] ;
assign n368 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n369 =  ( n368 ) == ( 16'd2 )  ;
assign n370 = aes_counter[23:16] ;
assign n371 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n372 =  ( n371 ) == ( 16'd1 )  ;
assign n373 = aes_counter[15:8] ;
assign n374 = aes_counter[7:0] ;
assign n375 =  ( n372 ) ? ( n373 ) : ( n374 ) ;
assign n376 =  ( n369 ) ? ( n370 ) : ( n375 ) ;
assign n377 =  ( n366 ) ? ( n367 ) : ( n376 ) ;
assign n378 =  ( n363 ) ? ( n364 ) : ( n377 ) ;
assign n379 =  ( n360 ) ? ( n361 ) : ( n378 ) ;
assign n380 =  ( n357 ) ? ( n358 ) : ( n379 ) ;
assign n381 =  ( n354 ) ? ( n355 ) : ( n380 ) ;
assign n382 =  ( n351 ) ? ( n352 ) : ( n381 ) ;
assign n383 =  ( n348 ) ? ( n349 ) : ( n382 ) ;
assign n384 =  ( n345 ) ? ( n346 ) : ( n383 ) ;
assign n385 =  ( n342 ) ? ( n343 ) : ( n384 ) ;
assign n386 =  ( n339 ) ? ( n340 ) : ( n385 ) ;
assign n387 =  ( n336 ) ? ( n337 ) : ( n386 ) ;
assign n388 =  ( n333 ) ? ( n334 ) : ( n387 ) ;
assign n389 =  ( n330 ) ? ( n331 ) : ( n388 ) ;
assign n390 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n391 =  ( n390 ) == ( 16'd15 )  ;
assign n392 = aes_counter[127:120] ;
assign n393 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n394 =  ( n393 ) == ( 16'd14 )  ;
assign n395 = aes_counter[119:112] ;
assign n396 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n397 =  ( n396 ) == ( 16'd13 )  ;
assign n398 = aes_counter[111:104] ;
assign n399 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n400 =  ( n399 ) == ( 16'd12 )  ;
assign n401 = aes_counter[103:96] ;
assign n402 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n403 =  ( n402 ) == ( 16'd11 )  ;
assign n404 = aes_counter[95:88] ;
assign n405 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n406 =  ( n405 ) == ( 16'd10 )  ;
assign n407 = aes_counter[87:80] ;
assign n408 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n409 =  ( n408 ) == ( 16'd9 )  ;
assign n410 = aes_counter[79:72] ;
assign n411 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n412 =  ( n411 ) == ( 16'd8 )  ;
assign n413 = aes_counter[71:64] ;
assign n414 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n415 =  ( n414 ) == ( 16'd7 )  ;
assign n416 = aes_counter[63:56] ;
assign n417 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n418 =  ( n417 ) == ( 16'd6 )  ;
assign n419 = aes_counter[55:48] ;
assign n420 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n421 =  ( n420 ) == ( 16'd5 )  ;
assign n422 = aes_counter[47:40] ;
assign n423 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n424 =  ( n423 ) == ( 16'd4 )  ;
assign n425 = aes_counter[39:32] ;
assign n426 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n427 =  ( n426 ) == ( 16'd3 )  ;
assign n428 = aes_counter[31:24] ;
assign n429 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n430 =  ( n429 ) == ( 16'd2 )  ;
assign n431 = aes_counter[23:16] ;
assign n432 =  ( cmdaddr ) - ( 16'd65296 )  ;
assign n433 =  ( n432 ) == ( 16'd1 )  ;
assign n434 = aes_counter[15:8] ;
assign n435 = aes_counter[7:0] ;
assign n436 =  ( n433 ) ? ( n434 ) : ( n435 ) ;
assign n437 =  ( n430 ) ? ( n431 ) : ( n436 ) ;
assign n438 =  ( n427 ) ? ( n428 ) : ( n437 ) ;
assign n439 =  ( n424 ) ? ( n425 ) : ( n438 ) ;
assign n440 =  ( n421 ) ? ( n422 ) : ( n439 ) ;
assign n441 =  ( n418 ) ? ( n419 ) : ( n440 ) ;
assign n442 =  ( n415 ) ? ( n416 ) : ( n441 ) ;
assign n443 =  ( n412 ) ? ( n413 ) : ( n442 ) ;
assign n444 =  ( n409 ) ? ( n410 ) : ( n443 ) ;
assign n445 =  ( n406 ) ? ( n407 ) : ( n444 ) ;
assign n446 =  ( n403 ) ? ( n404 ) : ( n445 ) ;
assign n447 =  ( n400 ) ? ( n401 ) : ( n446 ) ;
assign n448 =  ( n397 ) ? ( n398 ) : ( n447 ) ;
assign n449 =  ( n394 ) ? ( n395 ) : ( n448 ) ;
assign n450 =  ( n391 ) ? ( n392 ) : ( n449 ) ;
always @(posedge clk) begin
   if(rst) begin
   end
   else if(__ILA_AES_valid__) begin
       if ( __ILA_AES_decode_of_START_ENCRYPT__ && __ILA_AES_grant__[1] ) begin
           aes_status <= n74;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_status <= n77;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_address <= n85;
       end else if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_address <= aes_address;
       end else if ( __ILA_AES_decode_of_WRITE_COUNTER__ && __ILA_AES_grant__[9] ) begin
           aes_address <= aes_address;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           aes_length <= aes_length;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_length <= n95;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_length <= aes_length;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_counter <= aes_counter;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_counter <= aes_counter;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_counter <= aes_counter;
       end else if ( __ILA_AES_decode_of_WRITE_COUNTER__ && __ILA_AES_grant__[9] ) begin
           aes_counter <= n177;
       end
       if ( __ILA_AES_decode_of_WRITE_ADDRESS__ && __ILA_AES_grant__[0] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_WRITE_LENGTH__ && __ILA_AES_grant__[7] ) begin
           aes_key <= aes_key;
       end else if ( __ILA_AES_decode_of_WRITE_KEY__ && __ILA_AES_grant__[8] ) begin
           aes_key <= n257;
       end else if ( __ILA_AES_decode_of_WRITE_COUNTER__ && __ILA_AES_grant__[9] ) begin
           aes_key <= aes_key;
       end
       if ( __ILA_AES_decode_of_READ_LENGTH__ && __ILA_AES_grant__[2] ) begin
           outdata <= n262;
       end else if ( __ILA_AES_decode_of_READ_ADDRESS__ && __ILA_AES_grant__[3] ) begin
           outdata <= n267;
       end else if ( __ILA_AES_decode_of_READ_KEY__ && __ILA_AES_grant__[4] ) begin
           outdata <= n328;
       end else if ( __ILA_AES_decode_of_READ_COUNTER__ && __ILA_AES_grant__[5] ) begin
           outdata <= n389;
       end else if ( __ILA_AES_decode_of_GET_STATUS__ && __ILA_AES_grant__[6] ) begin
           outdata <= n450;
       end
   end
end
endmodule
